VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_asap7_64x256_1rw
  FOREIGN sram_asap7_64x256_1rw 0 0 ;
  SYMMETRY X Y ;
  SIZE 16.720 BY 33.600 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.288 0.024 0.312 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.528 0.024 0.552 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.768 0.024 0.792 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.008 0.024 1.032 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.248 0.024 1.272 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.488 0.024 1.512 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.728 0.024 1.752 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.968 0.024 1.992 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.208 0.024 2.232 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.448 0.024 2.472 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.688 0.024 2.712 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.928 0.024 2.952 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.168 0.024 3.192 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.408 0.024 3.432 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.648 0.024 3.672 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.888 0.024 3.912 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.128 0.024 4.152 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.368 0.024 4.392 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.608 0.024 4.632 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.848 0.024 4.872 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.088 0.024 5.112 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.328 0.024 5.352 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.568 0.024 5.592 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.808 0.024 5.832 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.048 0.024 6.072 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.288 0.024 6.312 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.528 0.024 6.552 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.768 0.024 6.792 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.008 0.024 7.032 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.248 0.024 7.272 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.488 0.024 7.512 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.728 0.024 7.752 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.968 0.024 7.992 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.208 0.024 8.232 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.448 0.024 8.472 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.688 0.024 8.712 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.928 0.024 8.952 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.168 0.024 9.192 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.408 0.024 9.432 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.648 0.024 9.672 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.888 0.024 9.912 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.128 0.024 10.152 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.368 0.024 10.392 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.608 0.024 10.632 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.848 0.024 10.872 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.088 0.024 11.112 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.328 0.024 11.352 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.568 0.024 11.592 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.808 0.024 11.832 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.048 0.024 12.072 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.288 0.024 12.312 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.528 0.024 12.552 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.768 0.024 12.792 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.008 0.024 13.032 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.248 0.024 13.272 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.488 0.024 13.512 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.728 0.024 13.752 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.968 0.024 13.992 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.208 0.024 14.232 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.448 0.024 14.472 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.688 0.024 14.712 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.928 0.024 14.952 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.168 0.024 15.192 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.216 0.024 15.240 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.456 0.024 15.480 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.696 0.024 15.720 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.936 0.024 15.960 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.176 0.024 16.200 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.416 0.024 16.440 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.656 0.024 16.680 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.896 0.024 16.920 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.136 0.024 17.160 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.376 0.024 17.400 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.616 0.024 17.640 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.856 0.024 17.880 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.096 0.024 18.120 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.336 0.024 18.360 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.576 0.024 18.600 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.816 0.024 18.840 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.056 0.024 19.080 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.296 0.024 19.320 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.536 0.024 19.560 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.776 0.024 19.800 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.016 0.024 20.040 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.256 0.024 20.280 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.496 0.024 20.520 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.736 0.024 20.760 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.976 0.024 21.000 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.216 0.024 21.240 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.456 0.024 21.480 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.696 0.024 21.720 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.936 0.024 21.960 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.176 0.024 22.200 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.416 0.024 22.440 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.656 0.024 22.680 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.896 0.024 22.920 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.136 0.024 23.160 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.376 0.024 23.400 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.616 0.024 23.640 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.856 0.024 23.880 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.096 0.024 24.120 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.336 0.024 24.360 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.576 0.024 24.600 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.816 0.024 24.840 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.056 0.024 25.080 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.296 0.024 25.320 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.536 0.024 25.560 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.776 0.024 25.800 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.016 0.024 26.040 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.256 0.024 26.280 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.496 0.024 26.520 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.736 0.024 26.760 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.976 0.024 27.000 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.216 0.024 27.240 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.456 0.024 27.480 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.696 0.024 27.720 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.936 0.024 27.960 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.176 0.024 28.200 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.416 0.024 28.440 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.656 0.024 28.680 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.896 0.024 28.920 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.136 0.024 29.160 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.376 0.024 29.400 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.616 0.024 29.640 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.856 0.024 29.880 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.096 0.024 30.120 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.336 0.024 30.360 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.384 0.024 30.408 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.624 0.024 30.648 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.864 0.024 30.888 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.104 0.024 31.128 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.344 0.024 31.368 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.584 0.024 31.608 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.824 0.024 31.848 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.064 0.024 32.088 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.112 0.024 32.136 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.352 0.024 32.376 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.592 0.024 32.616 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 16.672 0.096 ;
      RECT 0.048 0.768 16.672 0.864 ;
      RECT 0.048 1.536 16.672 1.632 ;
      RECT 0.048 2.304 16.672 2.400 ;
      RECT 0.048 3.072 16.672 3.168 ;
      RECT 0.048 3.840 16.672 3.936 ;
      RECT 0.048 4.608 16.672 4.704 ;
      RECT 0.048 5.376 16.672 5.472 ;
      RECT 0.048 6.144 16.672 6.240 ;
      RECT 0.048 6.912 16.672 7.008 ;
      RECT 0.048 7.680 16.672 7.776 ;
      RECT 0.048 8.448 16.672 8.544 ;
      RECT 0.048 9.216 16.672 9.312 ;
      RECT 0.048 9.984 16.672 10.080 ;
      RECT 0.048 10.752 16.672 10.848 ;
      RECT 0.048 11.520 16.672 11.616 ;
      RECT 0.048 12.288 16.672 12.384 ;
      RECT 0.048 13.056 16.672 13.152 ;
      RECT 0.048 13.824 16.672 13.920 ;
      RECT 0.048 14.592 16.672 14.688 ;
      RECT 0.048 15.360 16.672 15.456 ;
      RECT 0.048 16.128 16.672 16.224 ;
      RECT 0.048 16.896 16.672 16.992 ;
      RECT 0.048 17.664 16.672 17.760 ;
      RECT 0.048 18.432 16.672 18.528 ;
      RECT 0.048 19.200 16.672 19.296 ;
      RECT 0.048 19.968 16.672 20.064 ;
      RECT 0.048 20.736 16.672 20.832 ;
      RECT 0.048 21.504 16.672 21.600 ;
      RECT 0.048 22.272 16.672 22.368 ;
      RECT 0.048 23.040 16.672 23.136 ;
      RECT 0.048 23.808 16.672 23.904 ;
      RECT 0.048 24.576 16.672 24.672 ;
      RECT 0.048 25.344 16.672 25.440 ;
      RECT 0.048 26.112 16.672 26.208 ;
      RECT 0.048 26.880 16.672 26.976 ;
      RECT 0.048 27.648 16.672 27.744 ;
      RECT 0.048 28.416 16.672 28.512 ;
      RECT 0.048 29.184 16.672 29.280 ;
      RECT 0.048 29.952 16.672 30.048 ;
      RECT 0.048 30.720 16.672 30.816 ;
      RECT 0.048 31.488 16.672 31.584 ;
      RECT 0.048 32.256 16.672 32.352 ;
      RECT 0.048 33.024 16.672 33.120 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 16.672 0.480 ;
      RECT 0.048 1.152 16.672 1.248 ;
      RECT 0.048 1.920 16.672 2.016 ;
      RECT 0.048 2.688 16.672 2.784 ;
      RECT 0.048 3.456 16.672 3.552 ;
      RECT 0.048 4.224 16.672 4.320 ;
      RECT 0.048 4.992 16.672 5.088 ;
      RECT 0.048 5.760 16.672 5.856 ;
      RECT 0.048 6.528 16.672 6.624 ;
      RECT 0.048 7.296 16.672 7.392 ;
      RECT 0.048 8.064 16.672 8.160 ;
      RECT 0.048 8.832 16.672 8.928 ;
      RECT 0.048 9.600 16.672 9.696 ;
      RECT 0.048 10.368 16.672 10.464 ;
      RECT 0.048 11.136 16.672 11.232 ;
      RECT 0.048 11.904 16.672 12.000 ;
      RECT 0.048 12.672 16.672 12.768 ;
      RECT 0.048 13.440 16.672 13.536 ;
      RECT 0.048 14.208 16.672 14.304 ;
      RECT 0.048 14.976 16.672 15.072 ;
      RECT 0.048 15.744 16.672 15.840 ;
      RECT 0.048 16.512 16.672 16.608 ;
      RECT 0.048 17.280 16.672 17.376 ;
      RECT 0.048 18.048 16.672 18.144 ;
      RECT 0.048 18.816 16.672 18.912 ;
      RECT 0.048 19.584 16.672 19.680 ;
      RECT 0.048 20.352 16.672 20.448 ;
      RECT 0.048 21.120 16.672 21.216 ;
      RECT 0.048 21.888 16.672 21.984 ;
      RECT 0.048 22.656 16.672 22.752 ;
      RECT 0.048 23.424 16.672 23.520 ;
      RECT 0.048 24.192 16.672 24.288 ;
      RECT 0.048 24.960 16.672 25.056 ;
      RECT 0.048 25.728 16.672 25.824 ;
      RECT 0.048 26.496 16.672 26.592 ;
      RECT 0.048 27.264 16.672 27.360 ;
      RECT 0.048 28.032 16.672 28.128 ;
      RECT 0.048 28.800 16.672 28.896 ;
      RECT 0.048 29.568 16.672 29.664 ;
      RECT 0.048 30.336 16.672 30.432 ;
      RECT 0.048 31.104 16.672 31.200 ;
      RECT 0.048 31.872 16.672 31.968 ;
      RECT 0.048 32.640 16.672 32.736 ;
      RECT 0.048 33.408 16.672 33.504 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 16.720 33.600 ;
    LAYER M2 ;
    RECT 0 0 16.720 33.600 ;
    LAYER M3 ;
    RECT 0 0 16.720 33.600 ;
    LAYER M4 ;
    RECT 0.024 0 0.048 33.600 ;
    RECT 16.672 0 16.720 33.600 ;
    RECT 0.048 0.000 16.672 0.000 ;
    RECT 0.048 0.096 16.672 0.384 ;
    RECT 0.048 0.480 16.672 0.768 ;
    RECT 0.048 0.864 16.672 1.152 ;
    RECT 0.048 1.248 16.672 1.536 ;
    RECT 0.048 1.632 16.672 1.920 ;
    RECT 0.048 2.016 16.672 2.304 ;
    RECT 0.048 2.400 16.672 2.688 ;
    RECT 0.048 2.784 16.672 3.072 ;
    RECT 0.048 3.168 16.672 3.456 ;
    RECT 0.048 3.552 16.672 3.840 ;
    RECT 0.048 3.936 16.672 4.224 ;
    RECT 0.048 4.320 16.672 4.608 ;
    RECT 0.048 4.704 16.672 4.992 ;
    RECT 0.048 5.088 16.672 5.376 ;
    RECT 0.048 5.472 16.672 5.760 ;
    RECT 0.048 5.856 16.672 6.144 ;
    RECT 0.048 6.240 16.672 6.528 ;
    RECT 0.048 6.624 16.672 6.912 ;
    RECT 0.048 7.008 16.672 7.296 ;
    RECT 0.048 7.392 16.672 7.680 ;
    RECT 0.048 7.776 16.672 8.064 ;
    RECT 0.048 8.160 16.672 8.448 ;
    RECT 0.048 8.544 16.672 8.832 ;
    RECT 0.048 8.928 16.672 9.216 ;
    RECT 0.048 9.312 16.672 9.600 ;
    RECT 0.048 9.696 16.672 9.984 ;
    RECT 0.048 10.080 16.672 10.368 ;
    RECT 0.048 10.464 16.672 10.752 ;
    RECT 0.048 10.848 16.672 11.136 ;
    RECT 0.048 11.232 16.672 11.520 ;
    RECT 0.048 11.616 16.672 11.904 ;
    RECT 0.048 12.000 16.672 12.288 ;
    RECT 0.048 12.384 16.672 12.672 ;
    RECT 0.048 12.768 16.672 13.056 ;
    RECT 0.048 13.152 16.672 13.440 ;
    RECT 0.048 13.536 16.672 13.824 ;
    RECT 0.048 13.920 16.672 14.208 ;
    RECT 0.048 14.304 16.672 14.592 ;
    RECT 0.048 14.688 16.672 14.976 ;
    RECT 0.048 15.072 16.672 15.360 ;
    RECT 0.048 15.456 16.672 15.744 ;
    RECT 0.048 15.840 16.672 16.128 ;
    RECT 0.048 16.224 16.672 16.512 ;
    RECT 0.048 16.608 16.672 16.896 ;
    RECT 0.048 16.992 16.672 17.280 ;
    RECT 0.048 17.376 16.672 17.664 ;
    RECT 0.048 17.760 16.672 18.048 ;
    RECT 0.048 18.144 16.672 18.432 ;
    RECT 0.048 18.528 16.672 18.816 ;
    RECT 0.048 18.912 16.672 19.200 ;
    RECT 0.048 19.296 16.672 19.584 ;
    RECT 0.048 19.680 16.672 19.968 ;
    RECT 0.048 20.064 16.672 20.352 ;
    RECT 0.048 20.448 16.672 20.736 ;
    RECT 0.048 20.832 16.672 21.120 ;
    RECT 0.048 21.216 16.672 21.504 ;
    RECT 0.048 21.600 16.672 21.888 ;
    RECT 0.048 21.984 16.672 22.272 ;
    RECT 0.048 22.368 16.672 22.656 ;
    RECT 0.048 22.752 16.672 23.040 ;
    RECT 0.048 23.136 16.672 23.424 ;
    RECT 0.048 23.520 16.672 23.808 ;
    RECT 0.048 23.904 16.672 24.192 ;
    RECT 0.048 24.288 16.672 24.576 ;
    RECT 0.048 24.672 16.672 24.960 ;
    RECT 0.048 25.056 16.672 25.344 ;
    RECT 0.048 25.440 16.672 25.728 ;
    RECT 0.048 25.824 16.672 26.112 ;
    RECT 0.048 26.208 16.672 26.496 ;
    RECT 0.048 26.592 16.672 26.880 ;
    RECT 0.048 26.976 16.672 27.264 ;
    RECT 0.048 27.360 16.672 27.648 ;
    RECT 0.048 27.744 16.672 28.032 ;
    RECT 0.048 28.128 16.672 28.416 ;
    RECT 0.048 28.512 16.672 28.800 ;
    RECT 0.048 28.896 16.672 29.184 ;
    RECT 0.048 29.280 16.672 29.568 ;
    RECT 0.048 29.664 16.672 29.952 ;
    RECT 0.048 30.048 16.672 30.336 ;
    RECT 0.048 30.432 16.672 30.720 ;
    RECT 0.048 30.816 16.672 31.104 ;
    RECT 0.048 31.200 16.672 31.488 ;
    RECT 0.048 31.584 16.672 31.872 ;
    RECT 0.048 31.968 16.672 32.256 ;
    RECT 0.048 32.352 16.672 32.640 ;
    RECT 0.048 32.736 16.672 33.024 ;
    RECT 0.048 33.120 16.672 33.408 ;
    RECT 0.048 33.504 16.672 33.600 ;
    RECT 0 0.000 0.024 0.048 ;
    RECT 0 0.072 0.024 0.288 ;
    RECT 0 0.312 0.024 0.528 ;
    RECT 0 0.552 0.024 0.768 ;
    RECT 0 0.792 0.024 1.008 ;
    RECT 0 1.032 0.024 1.248 ;
    RECT 0 1.272 0.024 1.488 ;
    RECT 0 1.512 0.024 1.728 ;
    RECT 0 1.752 0.024 1.968 ;
    RECT 0 1.992 0.024 2.208 ;
    RECT 0 2.232 0.024 2.448 ;
    RECT 0 2.472 0.024 2.688 ;
    RECT 0 2.712 0.024 2.928 ;
    RECT 0 2.952 0.024 3.168 ;
    RECT 0 3.192 0.024 3.408 ;
    RECT 0 3.432 0.024 3.648 ;
    RECT 0 3.672 0.024 3.888 ;
    RECT 0 3.912 0.024 4.128 ;
    RECT 0 4.152 0.024 4.368 ;
    RECT 0 4.392 0.024 4.608 ;
    RECT 0 4.632 0.024 4.848 ;
    RECT 0 4.872 0.024 5.088 ;
    RECT 0 5.112 0.024 5.328 ;
    RECT 0 5.352 0.024 5.568 ;
    RECT 0 5.592 0.024 5.808 ;
    RECT 0 5.832 0.024 6.048 ;
    RECT 0 6.072 0.024 6.288 ;
    RECT 0 6.312 0.024 6.528 ;
    RECT 0 6.552 0.024 6.768 ;
    RECT 0 6.792 0.024 7.008 ;
    RECT 0 7.032 0.024 7.248 ;
    RECT 0 7.272 0.024 7.488 ;
    RECT 0 7.512 0.024 7.728 ;
    RECT 0 7.752 0.024 7.968 ;
    RECT 0 7.992 0.024 8.208 ;
    RECT 0 8.232 0.024 8.448 ;
    RECT 0 8.472 0.024 8.688 ;
    RECT 0 8.712 0.024 8.928 ;
    RECT 0 8.952 0.024 9.168 ;
    RECT 0 9.192 0.024 9.408 ;
    RECT 0 9.432 0.024 9.648 ;
    RECT 0 9.672 0.024 9.888 ;
    RECT 0 9.912 0.024 10.128 ;
    RECT 0 10.152 0.024 10.368 ;
    RECT 0 10.392 0.024 10.608 ;
    RECT 0 10.632 0.024 10.848 ;
    RECT 0 10.872 0.024 11.088 ;
    RECT 0 11.112 0.024 11.328 ;
    RECT 0 11.352 0.024 11.568 ;
    RECT 0 11.592 0.024 11.808 ;
    RECT 0 11.832 0.024 12.048 ;
    RECT 0 12.072 0.024 12.288 ;
    RECT 0 12.312 0.024 12.528 ;
    RECT 0 12.552 0.024 12.768 ;
    RECT 0 12.792 0.024 13.008 ;
    RECT 0 13.032 0.024 13.248 ;
    RECT 0 13.272 0.024 13.488 ;
    RECT 0 13.512 0.024 13.728 ;
    RECT 0 13.752 0.024 13.968 ;
    RECT 0 13.992 0.024 14.208 ;
    RECT 0 14.232 0.024 14.448 ;
    RECT 0 14.472 0.024 14.688 ;
    RECT 0 14.712 0.024 14.928 ;
    RECT 0 14.952 0.024 15.168 ;
    RECT 0 15.192 0.024 15.216 ;
    RECT 0 15.240 0.024 15.456 ;
    RECT 0 15.480 0.024 15.696 ;
    RECT 0 15.720 0.024 15.936 ;
    RECT 0 15.960 0.024 16.176 ;
    RECT 0 16.200 0.024 16.416 ;
    RECT 0 16.440 0.024 16.656 ;
    RECT 0 16.680 0.024 16.896 ;
    RECT 0 16.920 0.024 17.136 ;
    RECT 0 17.160 0.024 17.376 ;
    RECT 0 17.400 0.024 17.616 ;
    RECT 0 17.640 0.024 17.856 ;
    RECT 0 17.880 0.024 18.096 ;
    RECT 0 18.120 0.024 18.336 ;
    RECT 0 18.360 0.024 18.576 ;
    RECT 0 18.600 0.024 18.816 ;
    RECT 0 18.840 0.024 19.056 ;
    RECT 0 19.080 0.024 19.296 ;
    RECT 0 19.320 0.024 19.536 ;
    RECT 0 19.560 0.024 19.776 ;
    RECT 0 19.800 0.024 20.016 ;
    RECT 0 20.040 0.024 20.256 ;
    RECT 0 20.280 0.024 20.496 ;
    RECT 0 20.520 0.024 20.736 ;
    RECT 0 20.760 0.024 20.976 ;
    RECT 0 21.000 0.024 21.216 ;
    RECT 0 21.240 0.024 21.456 ;
    RECT 0 21.480 0.024 21.696 ;
    RECT 0 21.720 0.024 21.936 ;
    RECT 0 21.960 0.024 22.176 ;
    RECT 0 22.200 0.024 22.416 ;
    RECT 0 22.440 0.024 22.656 ;
    RECT 0 22.680 0.024 22.896 ;
    RECT 0 22.920 0.024 23.136 ;
    RECT 0 23.160 0.024 23.376 ;
    RECT 0 23.400 0.024 23.616 ;
    RECT 0 23.640 0.024 23.856 ;
    RECT 0 23.880 0.024 24.096 ;
    RECT 0 24.120 0.024 24.336 ;
    RECT 0 24.360 0.024 24.576 ;
    RECT 0 24.600 0.024 24.816 ;
    RECT 0 24.840 0.024 25.056 ;
    RECT 0 25.080 0.024 25.296 ;
    RECT 0 25.320 0.024 25.536 ;
    RECT 0 25.560 0.024 25.776 ;
    RECT 0 25.800 0.024 26.016 ;
    RECT 0 26.040 0.024 26.256 ;
    RECT 0 26.280 0.024 26.496 ;
    RECT 0 26.520 0.024 26.736 ;
    RECT 0 26.760 0.024 26.976 ;
    RECT 0 27.000 0.024 27.216 ;
    RECT 0 27.240 0.024 27.456 ;
    RECT 0 27.480 0.024 27.696 ;
    RECT 0 27.720 0.024 27.936 ;
    RECT 0 27.960 0.024 28.176 ;
    RECT 0 28.200 0.024 28.416 ;
    RECT 0 28.440 0.024 28.656 ;
    RECT 0 28.680 0.024 28.896 ;
    RECT 0 28.920 0.024 29.136 ;
    RECT 0 29.160 0.024 29.376 ;
    RECT 0 29.400 0.024 29.616 ;
    RECT 0 29.640 0.024 29.856 ;
    RECT 0 29.880 0.024 30.096 ;
    RECT 0 30.120 0.024 30.336 ;
    RECT 0 30.360 0.024 30.384 ;
    RECT 0 30.408 0.024 30.624 ;
    RECT 0 30.648 0.024 30.864 ;
    RECT 0 30.888 0.024 31.104 ;
    RECT 0 31.128 0.024 31.344 ;
    RECT 0 31.368 0.024 31.584 ;
    RECT 0 31.608 0.024 31.824 ;
    RECT 0 31.848 0.024 32.064 ;
    RECT 0 32.088 0.024 32.304 ;
    RECT 0 32.328 0.024 32.544 ;
    RECT 0 32.568 0.024 32.784 ;
    RECT 0 32.808 0.024 33.024 ;
    RECT 0 33.048 0.024 33.264 ;
    RECT 0 33.288 0.024 33.504 ;
    RECT 0 33.528 0.024 33.600 ;
  END
END sram_asap7_64x256_1rw

END LIBRARY
