VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_asap7_32x256_1rw
  FOREIGN sram_asap7_32x256_1rw 0 0 ;
  SYMMETRY X Y ;
  SIZE 16.720 BY 16.800 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.240 0.024 0.264 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.432 0.024 0.456 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.624 0.024 0.648 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.816 0.024 0.840 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.008 0.024 1.032 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.200 0.024 1.224 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.392 0.024 1.416 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.584 0.024 1.608 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.776 0.024 1.800 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.968 0.024 1.992 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.160 0.024 2.184 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.352 0.024 2.376 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.544 0.024 2.568 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.736 0.024 2.760 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.928 0.024 2.952 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.120 0.024 3.144 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.312 0.024 3.336 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.504 0.024 3.528 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.696 0.024 3.720 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.888 0.024 3.912 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.080 0.024 4.104 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.272 0.024 4.296 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.464 0.024 4.488 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.656 0.024 4.680 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.848 0.024 4.872 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.040 0.024 5.064 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.232 0.024 5.256 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.424 0.024 5.448 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.616 0.024 5.640 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.808 0.024 5.832 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.000 0.024 6.024 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.576 0.024 6.600 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.768 0.024 6.792 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.960 0.024 6.984 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.152 0.024 7.176 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.344 0.024 7.368 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.536 0.024 7.560 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.728 0.024 7.752 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.920 0.024 7.944 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.112 0.024 8.136 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.304 0.024 8.328 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.496 0.024 8.520 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.688 0.024 8.712 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.880 0.024 8.904 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.072 0.024 9.096 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.264 0.024 9.288 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.456 0.024 9.480 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.648 0.024 9.672 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.840 0.024 9.864 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.032 0.024 10.056 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.224 0.024 10.248 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.416 0.024 10.440 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.608 0.024 10.632 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.800 0.024 10.824 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.992 0.024 11.016 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.184 0.024 11.208 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.376 0.024 11.400 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.568 0.024 11.592 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.760 0.024 11.784 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.952 0.024 11.976 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.144 0.024 12.168 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.336 0.024 12.360 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.528 0.024 12.552 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.104 0.024 13.128 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.296 0.024 13.320 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.488 0.024 13.512 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.680 0.024 13.704 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.872 0.024 13.896 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.064 0.024 14.088 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.256 0.024 14.280 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.448 0.024 14.472 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.024 0.024 15.048 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.216 0.024 15.240 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.408 0.024 15.432 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 16.672 0.096 ;
      RECT 0.048 0.768 16.672 0.864 ;
      RECT 0.048 1.536 16.672 1.632 ;
      RECT 0.048 2.304 16.672 2.400 ;
      RECT 0.048 3.072 16.672 3.168 ;
      RECT 0.048 3.840 16.672 3.936 ;
      RECT 0.048 4.608 16.672 4.704 ;
      RECT 0.048 5.376 16.672 5.472 ;
      RECT 0.048 6.144 16.672 6.240 ;
      RECT 0.048 6.912 16.672 7.008 ;
      RECT 0.048 7.680 16.672 7.776 ;
      RECT 0.048 8.448 16.672 8.544 ;
      RECT 0.048 9.216 16.672 9.312 ;
      RECT 0.048 9.984 16.672 10.080 ;
      RECT 0.048 10.752 16.672 10.848 ;
      RECT 0.048 11.520 16.672 11.616 ;
      RECT 0.048 12.288 16.672 12.384 ;
      RECT 0.048 13.056 16.672 13.152 ;
      RECT 0.048 13.824 16.672 13.920 ;
      RECT 0.048 14.592 16.672 14.688 ;
      RECT 0.048 15.360 16.672 15.456 ;
      RECT 0.048 16.128 16.672 16.224 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 16.672 0.480 ;
      RECT 0.048 1.152 16.672 1.248 ;
      RECT 0.048 1.920 16.672 2.016 ;
      RECT 0.048 2.688 16.672 2.784 ;
      RECT 0.048 3.456 16.672 3.552 ;
      RECT 0.048 4.224 16.672 4.320 ;
      RECT 0.048 4.992 16.672 5.088 ;
      RECT 0.048 5.760 16.672 5.856 ;
      RECT 0.048 6.528 16.672 6.624 ;
      RECT 0.048 7.296 16.672 7.392 ;
      RECT 0.048 8.064 16.672 8.160 ;
      RECT 0.048 8.832 16.672 8.928 ;
      RECT 0.048 9.600 16.672 9.696 ;
      RECT 0.048 10.368 16.672 10.464 ;
      RECT 0.048 11.136 16.672 11.232 ;
      RECT 0.048 11.904 16.672 12.000 ;
      RECT 0.048 12.672 16.672 12.768 ;
      RECT 0.048 13.440 16.672 13.536 ;
      RECT 0.048 14.208 16.672 14.304 ;
      RECT 0.048 14.976 16.672 15.072 ;
      RECT 0.048 15.744 16.672 15.840 ;
      RECT 0.048 16.512 16.672 16.608 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 16.720 16.800 ;
    LAYER M2 ;
    RECT 0 0 16.720 16.800 ;
    LAYER M3 ;
    RECT 0 0 16.720 16.800 ;
    LAYER M4 ;
    RECT 0.024 0 0.048 16.800 ;
    RECT 16.672 0 16.720 16.800 ;
    RECT 0.048 0.000 16.672 0.000 ;
    RECT 0.048 0.096 16.672 0.384 ;
    RECT 0.048 0.480 16.672 0.768 ;
    RECT 0.048 0.864 16.672 1.152 ;
    RECT 0.048 1.248 16.672 1.536 ;
    RECT 0.048 1.632 16.672 1.920 ;
    RECT 0.048 2.016 16.672 2.304 ;
    RECT 0.048 2.400 16.672 2.688 ;
    RECT 0.048 2.784 16.672 3.072 ;
    RECT 0.048 3.168 16.672 3.456 ;
    RECT 0.048 3.552 16.672 3.840 ;
    RECT 0.048 3.936 16.672 4.224 ;
    RECT 0.048 4.320 16.672 4.608 ;
    RECT 0.048 4.704 16.672 4.992 ;
    RECT 0.048 5.088 16.672 5.376 ;
    RECT 0.048 5.472 16.672 5.760 ;
    RECT 0.048 5.856 16.672 6.144 ;
    RECT 0.048 6.240 16.672 6.528 ;
    RECT 0.048 6.624 16.672 6.912 ;
    RECT 0.048 7.008 16.672 7.296 ;
    RECT 0.048 7.392 16.672 7.680 ;
    RECT 0.048 7.776 16.672 8.064 ;
    RECT 0.048 8.160 16.672 8.448 ;
    RECT 0.048 8.544 16.672 8.832 ;
    RECT 0.048 8.928 16.672 9.216 ;
    RECT 0.048 9.312 16.672 9.600 ;
    RECT 0.048 9.696 16.672 9.984 ;
    RECT 0.048 10.080 16.672 10.368 ;
    RECT 0.048 10.464 16.672 10.752 ;
    RECT 0.048 10.848 16.672 11.136 ;
    RECT 0.048 11.232 16.672 11.520 ;
    RECT 0.048 11.616 16.672 11.904 ;
    RECT 0.048 12.000 16.672 12.288 ;
    RECT 0.048 12.384 16.672 12.672 ;
    RECT 0.048 12.768 16.672 13.056 ;
    RECT 0.048 13.152 16.672 13.440 ;
    RECT 0.048 13.536 16.672 13.824 ;
    RECT 0.048 13.920 16.672 14.208 ;
    RECT 0.048 14.304 16.672 14.592 ;
    RECT 0.048 14.688 16.672 14.976 ;
    RECT 0.048 15.072 16.672 15.360 ;
    RECT 0.048 15.456 16.672 15.744 ;
    RECT 0.048 15.840 16.672 16.128 ;
    RECT 0.048 16.224 16.672 16.512 ;
    RECT 0.048 16.608 16.672 16.800 ;
    RECT 0 0.000 0.024 0.048 ;
    RECT 0 0.072 0.024 0.240 ;
    RECT 0 0.264 0.024 0.432 ;
    RECT 0 0.456 0.024 0.624 ;
    RECT 0 0.648 0.024 0.816 ;
    RECT 0 0.840 0.024 1.008 ;
    RECT 0 1.032 0.024 1.200 ;
    RECT 0 1.224 0.024 1.392 ;
    RECT 0 1.416 0.024 1.584 ;
    RECT 0 1.608 0.024 1.776 ;
    RECT 0 1.800 0.024 1.968 ;
    RECT 0 1.992 0.024 2.160 ;
    RECT 0 2.184 0.024 2.352 ;
    RECT 0 2.376 0.024 2.544 ;
    RECT 0 2.568 0.024 2.736 ;
    RECT 0 2.760 0.024 2.928 ;
    RECT 0 2.952 0.024 3.120 ;
    RECT 0 3.144 0.024 3.312 ;
    RECT 0 3.336 0.024 3.504 ;
    RECT 0 3.528 0.024 3.696 ;
    RECT 0 3.720 0.024 3.888 ;
    RECT 0 3.912 0.024 4.080 ;
    RECT 0 4.104 0.024 4.272 ;
    RECT 0 4.296 0.024 4.464 ;
    RECT 0 4.488 0.024 4.656 ;
    RECT 0 4.680 0.024 4.848 ;
    RECT 0 4.872 0.024 5.040 ;
    RECT 0 5.064 0.024 5.232 ;
    RECT 0 5.256 0.024 5.424 ;
    RECT 0 5.448 0.024 5.616 ;
    RECT 0 5.640 0.024 5.808 ;
    RECT 0 5.832 0.024 6.000 ;
    RECT 0 6.024 0.024 6.576 ;
    RECT 0 6.600 0.024 6.768 ;
    RECT 0 6.792 0.024 6.960 ;
    RECT 0 6.984 0.024 7.152 ;
    RECT 0 7.176 0.024 7.344 ;
    RECT 0 7.368 0.024 7.536 ;
    RECT 0 7.560 0.024 7.728 ;
    RECT 0 7.752 0.024 7.920 ;
    RECT 0 7.944 0.024 8.112 ;
    RECT 0 8.136 0.024 8.304 ;
    RECT 0 8.328 0.024 8.496 ;
    RECT 0 8.520 0.024 8.688 ;
    RECT 0 8.712 0.024 8.880 ;
    RECT 0 8.904 0.024 9.072 ;
    RECT 0 9.096 0.024 9.264 ;
    RECT 0 9.288 0.024 9.456 ;
    RECT 0 9.480 0.024 9.648 ;
    RECT 0 9.672 0.024 9.840 ;
    RECT 0 9.864 0.024 10.032 ;
    RECT 0 10.056 0.024 10.224 ;
    RECT 0 10.248 0.024 10.416 ;
    RECT 0 10.440 0.024 10.608 ;
    RECT 0 10.632 0.024 10.800 ;
    RECT 0 10.824 0.024 10.992 ;
    RECT 0 11.016 0.024 11.184 ;
    RECT 0 11.208 0.024 11.376 ;
    RECT 0 11.400 0.024 11.568 ;
    RECT 0 11.592 0.024 11.760 ;
    RECT 0 11.784 0.024 11.952 ;
    RECT 0 11.976 0.024 12.144 ;
    RECT 0 12.168 0.024 12.336 ;
    RECT 0 12.360 0.024 12.528 ;
    RECT 0 12.552 0.024 13.104 ;
    RECT 0 13.128 0.024 13.296 ;
    RECT 0 13.320 0.024 13.488 ;
    RECT 0 13.512 0.024 13.680 ;
    RECT 0 13.704 0.024 13.872 ;
    RECT 0 13.896 0.024 14.064 ;
    RECT 0 14.088 0.024 14.256 ;
    RECT 0 14.280 0.024 14.448 ;
    RECT 0 14.472 0.024 14.640 ;
    RECT 0 14.664 0.024 14.832 ;
    RECT 0 14.856 0.024 15.024 ;
    RECT 0 15.048 0.024 15.216 ;
    RECT 0 15.240 0.024 15.408 ;
    RECT 0 15.432 0.024 15.600 ;
    RECT 0 15.624 0.024 15.792 ;
    RECT 0 15.816 0.024 15.984 ;
    RECT 0 16.008 0.024 16.176 ;
    RECT 0 16.200 0.024 16.368 ;
    RECT 0 16.392 0.024 16.560 ;
    RECT 0 16.584 0.024 16.752 ;
    RECT 0 16.776 0.024 16.800 ;
  END
END sram_asap7_32x256_1rw

END LIBRARY
