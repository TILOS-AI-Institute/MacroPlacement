VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_asap7_64x64_1rw
  FOREIGN sram_asap7_64x64_1rw 0 0 ;
  SYMMETRY X Y ;
  SIZE 8.360 BY 16.800 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.144 0.024 0.168 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.240 0.024 0.264 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.336 0.024 0.360 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.432 0.024 0.456 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.528 0.024 0.552 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.624 0.024 0.648 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.720 0.024 0.744 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.816 0.024 0.840 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.912 0.024 0.936 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.008 0.024 1.032 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.104 0.024 1.128 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.200 0.024 1.224 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.296 0.024 1.320 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.392 0.024 1.416 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.488 0.024 1.512 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.584 0.024 1.608 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.680 0.024 1.704 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.776 0.024 1.800 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.872 0.024 1.896 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.968 0.024 1.992 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.064 0.024 2.088 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.160 0.024 2.184 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.256 0.024 2.280 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.352 0.024 2.376 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.448 0.024 2.472 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.544 0.024 2.568 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.640 0.024 2.664 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.736 0.024 2.760 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.832 0.024 2.856 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.928 0.024 2.952 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.024 0.024 3.048 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.120 0.024 3.144 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.216 0.024 3.240 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.312 0.024 3.336 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.408 0.024 3.432 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.504 0.024 3.528 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.600 0.024 3.624 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.696 0.024 3.720 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.792 0.024 3.816 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.888 0.024 3.912 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.984 0.024 4.008 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.080 0.024 4.104 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.176 0.024 4.200 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.272 0.024 4.296 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.368 0.024 4.392 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.464 0.024 4.488 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.560 0.024 4.584 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.656 0.024 4.680 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.752 0.024 4.776 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.848 0.024 4.872 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.944 0.024 4.968 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.040 0.024 5.064 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.136 0.024 5.160 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.232 0.024 5.256 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.328 0.024 5.352 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.424 0.024 5.448 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.520 0.024 5.544 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.616 0.024 5.640 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.712 0.024 5.736 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.808 0.024 5.832 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.904 0.024 5.928 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.000 0.024 6.024 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.096 0.024 6.120 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.960 0.024 6.984 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.056 0.024 7.080 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.152 0.024 7.176 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.248 0.024 7.272 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.344 0.024 7.368 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.440 0.024 7.464 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.536 0.024 7.560 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.632 0.024 7.656 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.728 0.024 7.752 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.824 0.024 7.848 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.920 0.024 7.944 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.016 0.024 8.040 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.112 0.024 8.136 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.208 0.024 8.232 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.304 0.024 8.328 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.400 0.024 8.424 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.496 0.024 8.520 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.592 0.024 8.616 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.688 0.024 8.712 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.784 0.024 8.808 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.880 0.024 8.904 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.976 0.024 9.000 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.072 0.024 9.096 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.168 0.024 9.192 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.264 0.024 9.288 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.360 0.024 9.384 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.456 0.024 9.480 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.552 0.024 9.576 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.648 0.024 9.672 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.744 0.024 9.768 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.840 0.024 9.864 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.936 0.024 9.960 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.032 0.024 10.056 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.128 0.024 10.152 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.224 0.024 10.248 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.320 0.024 10.344 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.416 0.024 10.440 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.512 0.024 10.536 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.608 0.024 10.632 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.704 0.024 10.728 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.800 0.024 10.824 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.896 0.024 10.920 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.992 0.024 11.016 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.088 0.024 11.112 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.184 0.024 11.208 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.280 0.024 11.304 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.376 0.024 11.400 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.472 0.024 11.496 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.568 0.024 11.592 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.664 0.024 11.688 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.760 0.024 11.784 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.856 0.024 11.880 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.952 0.024 11.976 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.048 0.024 12.072 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.144 0.024 12.168 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.240 0.024 12.264 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.336 0.024 12.360 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.432 0.024 12.456 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.528 0.024 12.552 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.624 0.024 12.648 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.720 0.024 12.744 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.816 0.024 12.840 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.912 0.024 12.936 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.008 0.024 13.032 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.872 0.024 13.896 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.968 0.024 13.992 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.064 0.024 14.088 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.160 0.024 14.184 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.256 0.024 14.280 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.352 0.024 14.376 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.216 0.024 15.240 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.312 0.024 15.336 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.408 0.024 15.432 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 8.312 0.096 ;
      RECT 0.048 0.768 8.312 0.864 ;
      RECT 0.048 1.536 8.312 1.632 ;
      RECT 0.048 2.304 8.312 2.400 ;
      RECT 0.048 3.072 8.312 3.168 ;
      RECT 0.048 3.840 8.312 3.936 ;
      RECT 0.048 4.608 8.312 4.704 ;
      RECT 0.048 5.376 8.312 5.472 ;
      RECT 0.048 6.144 8.312 6.240 ;
      RECT 0.048 6.912 8.312 7.008 ;
      RECT 0.048 7.680 8.312 7.776 ;
      RECT 0.048 8.448 8.312 8.544 ;
      RECT 0.048 9.216 8.312 9.312 ;
      RECT 0.048 9.984 8.312 10.080 ;
      RECT 0.048 10.752 8.312 10.848 ;
      RECT 0.048 11.520 8.312 11.616 ;
      RECT 0.048 12.288 8.312 12.384 ;
      RECT 0.048 13.056 8.312 13.152 ;
      RECT 0.048 13.824 8.312 13.920 ;
      RECT 0.048 14.592 8.312 14.688 ;
      RECT 0.048 15.360 8.312 15.456 ;
      RECT 0.048 16.128 8.312 16.224 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 8.312 0.480 ;
      RECT 0.048 1.152 8.312 1.248 ;
      RECT 0.048 1.920 8.312 2.016 ;
      RECT 0.048 2.688 8.312 2.784 ;
      RECT 0.048 3.456 8.312 3.552 ;
      RECT 0.048 4.224 8.312 4.320 ;
      RECT 0.048 4.992 8.312 5.088 ;
      RECT 0.048 5.760 8.312 5.856 ;
      RECT 0.048 6.528 8.312 6.624 ;
      RECT 0.048 7.296 8.312 7.392 ;
      RECT 0.048 8.064 8.312 8.160 ;
      RECT 0.048 8.832 8.312 8.928 ;
      RECT 0.048 9.600 8.312 9.696 ;
      RECT 0.048 10.368 8.312 10.464 ;
      RECT 0.048 11.136 8.312 11.232 ;
      RECT 0.048 11.904 8.312 12.000 ;
      RECT 0.048 12.672 8.312 12.768 ;
      RECT 0.048 13.440 8.312 13.536 ;
      RECT 0.048 14.208 8.312 14.304 ;
      RECT 0.048 14.976 8.312 15.072 ;
      RECT 0.048 15.744 8.312 15.840 ;
      RECT 0.048 16.512 8.312 16.608 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 8.360 16.800 ;
    LAYER M2 ;
    RECT 0 0 8.360 16.800 ;
    LAYER M3 ;
    RECT 0 0 8.360 16.800 ;
    LAYER M4 ;
    RECT 0.024 0 0.048 16.800 ;
    RECT 8.312 0 8.360 16.800 ;
    RECT 0.048 0.000 8.312 0.000 ;
    RECT 0.048 0.096 8.312 0.384 ;
    RECT 0.048 0.480 8.312 0.768 ;
    RECT 0.048 0.864 8.312 1.152 ;
    RECT 0.048 1.248 8.312 1.536 ;
    RECT 0.048 1.632 8.312 1.920 ;
    RECT 0.048 2.016 8.312 2.304 ;
    RECT 0.048 2.400 8.312 2.688 ;
    RECT 0.048 2.784 8.312 3.072 ;
    RECT 0.048 3.168 8.312 3.456 ;
    RECT 0.048 3.552 8.312 3.840 ;
    RECT 0.048 3.936 8.312 4.224 ;
    RECT 0.048 4.320 8.312 4.608 ;
    RECT 0.048 4.704 8.312 4.992 ;
    RECT 0.048 5.088 8.312 5.376 ;
    RECT 0.048 5.472 8.312 5.760 ;
    RECT 0.048 5.856 8.312 6.144 ;
    RECT 0.048 6.240 8.312 6.528 ;
    RECT 0.048 6.624 8.312 6.912 ;
    RECT 0.048 7.008 8.312 7.296 ;
    RECT 0.048 7.392 8.312 7.680 ;
    RECT 0.048 7.776 8.312 8.064 ;
    RECT 0.048 8.160 8.312 8.448 ;
    RECT 0.048 8.544 8.312 8.832 ;
    RECT 0.048 8.928 8.312 9.216 ;
    RECT 0.048 9.312 8.312 9.600 ;
    RECT 0.048 9.696 8.312 9.984 ;
    RECT 0.048 10.080 8.312 10.368 ;
    RECT 0.048 10.464 8.312 10.752 ;
    RECT 0.048 10.848 8.312 11.136 ;
    RECT 0.048 11.232 8.312 11.520 ;
    RECT 0.048 11.616 8.312 11.904 ;
    RECT 0.048 12.000 8.312 12.288 ;
    RECT 0.048 12.384 8.312 12.672 ;
    RECT 0.048 12.768 8.312 13.056 ;
    RECT 0.048 13.152 8.312 13.440 ;
    RECT 0.048 13.536 8.312 13.824 ;
    RECT 0.048 13.920 8.312 14.208 ;
    RECT 0.048 14.304 8.312 14.592 ;
    RECT 0.048 14.688 8.312 14.976 ;
    RECT 0.048 15.072 8.312 15.360 ;
    RECT 0.048 15.456 8.312 15.744 ;
    RECT 0.048 15.840 8.312 16.128 ;
    RECT 0.048 16.224 8.312 16.512 ;
    RECT 0.048 16.608 8.312 16.800 ;
    RECT 0 0.000 0.024 0.048 ;
    RECT 0 0.072 0.024 0.144 ;
    RECT 0 0.168 0.024 0.240 ;
    RECT 0 0.264 0.024 0.336 ;
    RECT 0 0.360 0.024 0.432 ;
    RECT 0 0.456 0.024 0.528 ;
    RECT 0 0.552 0.024 0.624 ;
    RECT 0 0.648 0.024 0.720 ;
    RECT 0 0.744 0.024 0.816 ;
    RECT 0 0.840 0.024 0.912 ;
    RECT 0 0.936 0.024 1.008 ;
    RECT 0 1.032 0.024 1.104 ;
    RECT 0 1.128 0.024 1.200 ;
    RECT 0 1.224 0.024 1.296 ;
    RECT 0 1.320 0.024 1.392 ;
    RECT 0 1.416 0.024 1.488 ;
    RECT 0 1.512 0.024 1.584 ;
    RECT 0 1.608 0.024 1.680 ;
    RECT 0 1.704 0.024 1.776 ;
    RECT 0 1.800 0.024 1.872 ;
    RECT 0 1.896 0.024 1.968 ;
    RECT 0 1.992 0.024 2.064 ;
    RECT 0 2.088 0.024 2.160 ;
    RECT 0 2.184 0.024 2.256 ;
    RECT 0 2.280 0.024 2.352 ;
    RECT 0 2.376 0.024 2.448 ;
    RECT 0 2.472 0.024 2.544 ;
    RECT 0 2.568 0.024 2.640 ;
    RECT 0 2.664 0.024 2.736 ;
    RECT 0 2.760 0.024 2.832 ;
    RECT 0 2.856 0.024 2.928 ;
    RECT 0 2.952 0.024 3.024 ;
    RECT 0 3.048 0.024 3.120 ;
    RECT 0 3.144 0.024 3.216 ;
    RECT 0 3.240 0.024 3.312 ;
    RECT 0 3.336 0.024 3.408 ;
    RECT 0 3.432 0.024 3.504 ;
    RECT 0 3.528 0.024 3.600 ;
    RECT 0 3.624 0.024 3.696 ;
    RECT 0 3.720 0.024 3.792 ;
    RECT 0 3.816 0.024 3.888 ;
    RECT 0 3.912 0.024 3.984 ;
    RECT 0 4.008 0.024 4.080 ;
    RECT 0 4.104 0.024 4.176 ;
    RECT 0 4.200 0.024 4.272 ;
    RECT 0 4.296 0.024 4.368 ;
    RECT 0 4.392 0.024 4.464 ;
    RECT 0 4.488 0.024 4.560 ;
    RECT 0 4.584 0.024 4.656 ;
    RECT 0 4.680 0.024 4.752 ;
    RECT 0 4.776 0.024 4.848 ;
    RECT 0 4.872 0.024 4.944 ;
    RECT 0 4.968 0.024 5.040 ;
    RECT 0 5.064 0.024 5.136 ;
    RECT 0 5.160 0.024 5.232 ;
    RECT 0 5.256 0.024 5.328 ;
    RECT 0 5.352 0.024 5.424 ;
    RECT 0 5.448 0.024 5.520 ;
    RECT 0 5.544 0.024 5.616 ;
    RECT 0 5.640 0.024 5.712 ;
    RECT 0 5.736 0.024 5.808 ;
    RECT 0 5.832 0.024 5.904 ;
    RECT 0 5.928 0.024 6.000 ;
    RECT 0 6.024 0.024 6.096 ;
    RECT 0 6.120 0.024 6.960 ;
    RECT 0 6.984 0.024 7.056 ;
    RECT 0 7.080 0.024 7.152 ;
    RECT 0 7.176 0.024 7.248 ;
    RECT 0 7.272 0.024 7.344 ;
    RECT 0 7.368 0.024 7.440 ;
    RECT 0 7.464 0.024 7.536 ;
    RECT 0 7.560 0.024 7.632 ;
    RECT 0 7.656 0.024 7.728 ;
    RECT 0 7.752 0.024 7.824 ;
    RECT 0 7.848 0.024 7.920 ;
    RECT 0 7.944 0.024 8.016 ;
    RECT 0 8.040 0.024 8.112 ;
    RECT 0 8.136 0.024 8.208 ;
    RECT 0 8.232 0.024 8.304 ;
    RECT 0 8.328 0.024 8.400 ;
    RECT 0 8.424 0.024 8.496 ;
    RECT 0 8.520 0.024 8.592 ;
    RECT 0 8.616 0.024 8.688 ;
    RECT 0 8.712 0.024 8.784 ;
    RECT 0 8.808 0.024 8.880 ;
    RECT 0 8.904 0.024 8.976 ;
    RECT 0 9.000 0.024 9.072 ;
    RECT 0 9.096 0.024 9.168 ;
    RECT 0 9.192 0.024 9.264 ;
    RECT 0 9.288 0.024 9.360 ;
    RECT 0 9.384 0.024 9.456 ;
    RECT 0 9.480 0.024 9.552 ;
    RECT 0 9.576 0.024 9.648 ;
    RECT 0 9.672 0.024 9.744 ;
    RECT 0 9.768 0.024 9.840 ;
    RECT 0 9.864 0.024 9.936 ;
    RECT 0 9.960 0.024 10.032 ;
    RECT 0 10.056 0.024 10.128 ;
    RECT 0 10.152 0.024 10.224 ;
    RECT 0 10.248 0.024 10.320 ;
    RECT 0 10.344 0.024 10.416 ;
    RECT 0 10.440 0.024 10.512 ;
    RECT 0 10.536 0.024 10.608 ;
    RECT 0 10.632 0.024 10.704 ;
    RECT 0 10.728 0.024 10.800 ;
    RECT 0 10.824 0.024 10.896 ;
    RECT 0 10.920 0.024 10.992 ;
    RECT 0 11.016 0.024 11.088 ;
    RECT 0 11.112 0.024 11.184 ;
    RECT 0 11.208 0.024 11.280 ;
    RECT 0 11.304 0.024 11.376 ;
    RECT 0 11.400 0.024 11.472 ;
    RECT 0 11.496 0.024 11.568 ;
    RECT 0 11.592 0.024 11.664 ;
    RECT 0 11.688 0.024 11.760 ;
    RECT 0 11.784 0.024 11.856 ;
    RECT 0 11.880 0.024 11.952 ;
    RECT 0 11.976 0.024 12.048 ;
    RECT 0 12.072 0.024 12.144 ;
    RECT 0 12.168 0.024 12.240 ;
    RECT 0 12.264 0.024 12.336 ;
    RECT 0 12.360 0.024 12.432 ;
    RECT 0 12.456 0.024 12.528 ;
    RECT 0 12.552 0.024 12.624 ;
    RECT 0 12.648 0.024 12.720 ;
    RECT 0 12.744 0.024 12.816 ;
    RECT 0 12.840 0.024 12.912 ;
    RECT 0 12.936 0.024 13.008 ;
    RECT 0 13.032 0.024 13.872 ;
    RECT 0 13.896 0.024 13.968 ;
    RECT 0 13.992 0.024 14.064 ;
    RECT 0 14.088 0.024 14.160 ;
    RECT 0 14.184 0.024 14.256 ;
    RECT 0 14.280 0.024 14.352 ;
    RECT 0 14.376 0.024 14.448 ;
    RECT 0 14.472 0.024 14.544 ;
    RECT 0 14.568 0.024 14.640 ;
    RECT 0 14.664 0.024 14.736 ;
    RECT 0 14.760 0.024 14.832 ;
    RECT 0 14.856 0.024 14.928 ;
    RECT 0 14.952 0.024 15.024 ;
    RECT 0 15.048 0.024 15.120 ;
    RECT 0 15.144 0.024 15.216 ;
    RECT 0 15.240 0.024 15.312 ;
    RECT 0 15.336 0.024 15.408 ;
    RECT 0 15.432 0.024 15.504 ;
    RECT 0 15.528 0.024 15.600 ;
    RECT 0 15.624 0.024 15.696 ;
    RECT 0 15.720 0.024 15.792 ;
    RECT 0 15.816 0.024 15.888 ;
    RECT 0 15.912 0.024 15.984 ;
    RECT 0 16.008 0.024 16.080 ;
    RECT 0 16.104 0.024 16.176 ;
    RECT 0 16.200 0.024 16.272 ;
    RECT 0 16.296 0.024 16.368 ;
    RECT 0 16.392 0.024 16.464 ;
    RECT 0 16.488 0.024 16.560 ;
    RECT 0 16.584 0.024 16.656 ;
    RECT 0 16.680 0.024 16.752 ;
    RECT 0 16.776 0.024 16.848 ;
    RECT 0 16.872 0.024 16.944 ;
    RECT 0 16.968 0.024 17.040 ;
    RECT 0 17.064 0.024 17.136 ;
    RECT 0 17.160 0.024 17.232 ;
    RECT 0 17.256 0.024 17.328 ;
    RECT 0 17.352 0.024 17.424 ;
    RECT 0 17.448 0.024 17.520 ;
    RECT 0 17.544 0.024 17.616 ;
    RECT 0 17.640 0.024 17.712 ;
    RECT 0 17.736 0.024 17.808 ;
    RECT 0 17.832 0.024 17.904 ;
    RECT 0 17.928 0.024 18.000 ;
    RECT 0 18.024 0.024 18.096 ;
    RECT 0 18.120 0.024 18.192 ;
    RECT 0 18.216 0.024 18.288 ;
    RECT 0 18.312 0.024 18.384 ;
    RECT 0 18.408 0.024 18.480 ;
    RECT 0 18.504 0.024 18.576 ;
    RECT 0 18.600 0.024 18.672 ;
    RECT 0 18.696 0.024 18.768 ;
    RECT 0 18.792 0.024 18.864 ;
    RECT 0 18.888 0.024 18.960 ;
    RECT 0 18.984 0.024 19.056 ;
    RECT 0 19.080 0.024 19.152 ;
    RECT 0 19.176 0.024 19.248 ;
    RECT 0 19.272 0.024 19.344 ;
    RECT 0 19.368 0.024 19.440 ;
    RECT 0 19.464 0.024 19.536 ;
    RECT 0 19.560 0.024 19.632 ;
    RECT 0 19.656 0.024 19.728 ;
    RECT 0 19.752 0.024 19.824 ;
    RECT 0 19.848 0.024 19.920 ;
    RECT 0 19.944 0.024 20.784 ;
    RECT 0 20.808 0.024 20.880 ;
    RECT 0 20.904 0.024 20.976 ;
    RECT 0 21.000 0.024 21.072 ;
    RECT 0 21.096 0.024 21.168 ;
    RECT 0 21.192 0.024 21.264 ;
    RECT 0 21.288 0.024 22.128 ;
    RECT 0 22.152 0.024 22.224 ;
    RECT 0 22.248 0.024 22.320 ;
    RECT 0 22.344 0.024 16.800 ;
    LAYER OVERLAP ;
    RECT 0 0 8.360 16.800 ;
  END
END sram_asap7_64x64_1rw

END LIBRARY
