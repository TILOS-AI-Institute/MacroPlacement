VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

SITE FAKE_SITE_1H
  SIZE 0.057 BY 0.24 ;
  CLASS CORE ;
  SYMMETRY Y ;
END FAKE_SITE_1H

SITE FAKE_SITE_2H
  SIZE 0.057 BY 0.48 ;
  CLASS CORE ;
  SYMMETRY Y ;
END FAKE_SITE_2H

SITE FAKE_SITE_3H
  SIZE 0.057 BY 0.72 ;
  CLASS CORE ;
  SYMMETRY Y ;
END FAKE_SITE_3H

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.032 ;
  WIDTH 0.016 ;
  SPACING 0.016 ;
END M1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.016 ;
  WIDTH 0.016 ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.032 ;
  WIDTH 0.016 ;
  SPACING 0.016 ;
END M2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.016 ;
  WIDTH 0.016 ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.032 ;
  WIDTH 0.016 ;
  SPACING 0.016 ;
END M3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.016 ;
  WIDTH 0.016 ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.032 ;
  WIDTH 0.016 ;
  SPACING 0.016 ;
END M4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.016 ;
  WIDTH 0.016 ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.032 ;
  WIDTH 0.016 ;
  SPACING 0.016 ;
END M5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.016 ;
  WIDTH 0.016 ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.032 ;
  WIDTH 0.016 ;
  SPACING 0.016 ;
END M6

LAYER VIA6
  TYPE CUT ;
  SPACING 0.016 ;
  WIDTH 0.016 ;
END VIA6

MACRO SDFRPQD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.855 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END O1

END SDFRPQD1BWP240H8P57PDSVT


MACRO SDFRPQD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQD4BWP240H8P57PDSVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END SDFRPQD4BWP240H8P57PDSVT


MACRO CKLNQD12BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD12BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END CKLNQD12BWP240H8P57PDLVT


MACRO CKLNQOPTBBD12BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD12BWP240H8P57PDLVT 0 0 ;
  SIZE 1.083 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.24 0.5415 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.24 0.5415 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.24 0.5415 0.24 ;
    END
  END O1

END CKLNQOPTBBD12BWP240H8P57PDLVT


MACRO CKLNQD5BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD5BWP240H8P57PDLVT 0 0 ;
  SIZE 0.741 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END O1

END CKLNQD5BWP240H8P57PDLVT


MACRO CKLNQD6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END O1

END CKLNQD6BWP240H8P57PDLVT


MACRO CKLNQD6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END O1

END CKLNQD6BWP240H8P57PDSVT


MACRO CKLNQD14BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD14BWP240H8P57PDLVT 0 0 ;
  SIZE 1.083 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.24 0.5415 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.24 0.5415 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.24 0.5415 0.24 ;
    END
  END O1

END CKLNQD14BWP240H8P57PDLVT


MACRO CKLNQOPTBBD24BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD24BWP240H8P57PDLVT 0 0 ;
  SIZE 1.197 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.36 0.5985 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.36 0.5985 0.36 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.36 0.5985 0.36 ;
    END
  END O1

END CKLNQOPTBBD24BWP240H8P57PDLVT


MACRO CKLNQD16BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD16BWP240H8P57PDLVT 0 0 ;
  SIZE 0.855 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.36 0.4275 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.36 0.4275 0.36 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.36 0.4275 0.36 ;
    END
  END O1

END CKLNQD16BWP240H8P57PDLVT


MACRO CKLNQOPTBBD20BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD20BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.36 0.513 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.36 0.513 0.36 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.36 0.513 0.36 ;
    END
  END O1

END CKLNQOPTBBD20BWP240H8P57PDLVT


MACRO CKLNQD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END CKLNQD2BWP240H8P57PDSVT


MACRO CKLNQD24BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD24BWP240H8P57PDLVT 0 0 ;
  SIZE 1.197 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.36 0.5985 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.36 0.5985 0.36 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.36 0.5985 0.36 ;
    END
  END O1

END CKLNQD24BWP240H8P57PDLVT


MACRO CKLNQD20BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD20BWP240H8P57PDLVT 0 0 ;
  SIZE 0.969 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END O1

END CKLNQD20BWP240H8P57PDLVT


MACRO SDFSNQD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSNQD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END O1

END SDFSNQD1BWP240H8P57PDSVT


MACRO SDFRPQOPTQD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTQD2BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END SDFRPQOPTQD2BWP240H8P57PDLVT


MACRO SDFRPQD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END O1

END SDFRPQD2BWP240H8P57PDSVT


MACRO CKLNQD3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.24 0.3135 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.24 0.3135 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.24 0.3135 0.24 ;
    END
  END O1

END CKLNQD3BWP240H8P57PDLVT


MACRO CKLNQOPTBBD14BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD14BWP240H8P57PDLVT 0 0 ;
  SIZE 1.14 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END O1

END CKLNQOPTBBD14BWP240H8P57PDLVT


MACRO CKLNQOPTBBD8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD8BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END O1

END CKLNQOPTBBD8BWP240H8P57PDLVT


MACRO CKLNQOPTBBD10BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD10BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END CKLNQOPTBBD10BWP240H8P57PDLVT


MACRO CKLNQD10BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD10BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END O1

END CKLNQD10BWP240H8P57PDLVT


MACRO CKLNQOPTBBD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END O1

END CKLNQOPTBBD4BWP240H8P57PDLVT


MACRO CKLNQD3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.24 0.3135 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.24 0.3135 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.24 0.3135 0.24 ;
    END
  END O1

END CKLNQD3BWP240H8P57PDSVT


MACRO CKLNQD18BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD18BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END O1

END CKLNQD18BWP240H8P57PDLVT


MACRO CKLNQOPTBBD16BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQOPTBBD16BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END O1

END CKLNQOPTBBD16BWP240H8P57PDLVT


MACRO SDFRPQD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END O1

END SDFRPQD2BWP240H8P57PDLVT


MACRO SDFRPQOPTBBD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBBD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.969 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END O1

END SDFRPQOPTBBD1BWP240H8P57PDSVT


MACRO SDFRPQOPTBBD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBBD2BWP240H8P57PDSVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END SDFRPQOPTBBD2BWP240H8P57PDSVT


MACRO SDFRPQD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.855 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END O1

END SDFRPQD1BWP240H8P57PDLVT


MACRO CKLNQD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END CKLNQD2BWP240H8P57PDLVT


MACRO CKLNQD8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD8BWP240H8P57PDLVT 0 0 ;
  SIZE 0.855 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END O1

END CKLNQD8BWP240H8P57PDLVT


MACRO CKLNQD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKLNQD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END O1

END CKLNQD4BWP240H8P57PDLVT


MACRO SDFRPQOPTQD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTQD2BWP240H8P57PDSVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END SDFRPQOPTQD2BWP240H8P57PDSVT


MACRO SDFRPQD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQD4BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END SDFRPQD4BWP240H8P57PDLVT


MACRO SDFRPQOPTQD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTQD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.969 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END O1

END SDFRPQOPTQD1BWP240H8P57PDSVT


MACRO INVD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.171 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0855 0.12 0.0855 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0855 0.12 0.0855 0.12 ;
    END
  END O1

END INVD1BWP240H8P57PDSVT


MACRO INVD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END INVD2BWP240H8P57PDSVT


MACRO NR2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END NR2D1BWP240H8P57PDSVT


MACRO OAOI211D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OAOI211D1BWP240H8P57PDSVT


MACRO BUFFD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END BUFFD1BWP240H8P57PDSVT


MACRO BUFFD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END BUFFD2BWP240H8P57PDSVT


MACRO INVD3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END INVD3BWP240H8P57PDSVT


MACRO BUFFD5BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD5BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END BUFFD5BWP240H8P57PDSVT


MACRO BUFFD3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END BUFFD3BWP240H8P57PDSVT


MACRO XNR2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNR2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END XNR2D1BWP240H8P57PDSVT


MACRO ND2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END ND2D1BWP240H8P57PDSVT


MACRO OR2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END OR2D1BWP240H8P57PDSVT


MACRO OA21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OA21D1BWP240H8P57PDSVT


MACRO AOI21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END AOI21D1BWP240H8P57PDSVT


MACRO AN3D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN3D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AN3D2BWP240H8P57PDSVT


MACRO INR3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END INR3D1BWP240H8P57PDSVT


MACRO OAI211D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OAI211D1BWP240H8P57PDSVT


MACRO ND3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END ND3D1BWP240H8P57PDSVT


MACRO INR2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END INR2D1BWP240H8P57PDSVT


MACRO IAO21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAO21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END IAO21D1BWP240H8P57PDSVT


MACRO AOAI211D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOAI211D1BWP240H8P57PDSVT


MACRO AN2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END AN2D1BWP240H8P57PDSVT


MACRO AOI31D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOI31D1BWP240H8P57PDSVT


MACRO XOR2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END XOR2D1BWP240H8P57PDSVT


MACRO IND2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END IND2D1BWP240H8P57PDSVT


MACRO AOI22D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOI22D1BWP240H8P57PDSVT


MACRO AOI211D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOI211D1BWP240H8P57PDSVT


MACRO INR2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END INR2D2BWP240H8P57PDSVT


MACRO INR2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END INR2D4BWP240H8P57PDSVT


MACRO INR2D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END INR2D3BWP240H8P57PDSVT


MACRO OAI31D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OAI31D1BWP240H8P57PDSVT


MACRO OAI32D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OAI32D1BWP240H8P57PDSVT


MACRO OAI22D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OAI22D1BWP240H8P57PDSVT


MACRO OAI21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END OAI21D1BWP240H8P57PDSVT


MACRO AOI22D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOI22D1BWP240H8P57PDLVT


MACRO AO22D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AO22D1BWP240H8P57PDSVT


MACRO MOAI22D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MOAI22D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END MOAI22D2BWP240H8P57PDSVT


MACRO IOA21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END IOA21D1BWP240H8P57PDSVT


MACRO MOAI22D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MOAI22D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END MOAI22D2BWP240H8P57PDLVT


MACRO IAOI21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAOI21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END IAOI21D1BWP240H8P57PDSVT


MACRO XNR2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNR2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END XNR2D1BWP240H8P57PDLVT


MACRO AOI31D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOI31D1BWP240H8P57PDLVT


MACRO XNR2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNR2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END XNR2D2BWP240H8P57PDSVT


MACRO XNR2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNR2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END XNR2D2BWP240H8P57PDLVT


MACRO XOR2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END XOR2D2BWP240H8P57PDLVT


MACRO XOR2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END XOR2D1BWP240H8P57PDLVT


MACRO XOR2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END XOR2D2BWP240H8P57PDSVT


MACRO ND4D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END ND4D1BWP240H8P57PDSVT


MACRO ND4D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END ND4D1BWP240H8P57PDLVT


MACRO ND4SKFD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4SKFD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END ND4SKFD4BWP240H8P57PDLVT


MACRO ND4D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END O1

END ND4D3BWP240H8P57PDSVT


MACRO ND4D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END O1

END ND4D3BWP240H8P57PDLVT


MACRO BUFFD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END BUFFD4BWP240H8P57PDSVT


MACRO ND4D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END ND4D2BWP240H8P57PDSVT


MACRO NR4D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END NR4D1BWP240H8P57PDSVT


MACRO BUFFD5BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD5BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END BUFFD5BWP240H8P57PDLVT


MACRO INVD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END INVD4BWP240H8P57PDSVT


MACRO NR3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END NR3D1BWP240H8P57PDSVT


MACRO BUFFD8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD8BWP240H8P57PDSVT 0 0 ;
  SIZE 0.741 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END O1

END BUFFD8BWP240H8P57PDSVT


MACRO OR3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OR3D1BWP240H8P57PDSVT


MACRO NR2OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END NR2OPTPAD1BWP240H8P57PDSVT


MACRO ND2SKFD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2SKFD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END ND2SKFD4BWP240H8P57PDSVT


MACRO ND2SKFD3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2SKFD3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND2SKFD3BWP240H8P57PDSVT


MACRO BUFFD8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD8BWP240H8P57PDLVT 0 0 ;
  SIZE 0.741 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END O1

END BUFFD8BWP240H8P57PDLVT


MACRO INVD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END INVD2BWP240H8P57PDLVT


MACRO NR2D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END NR2D4BWP240H8P57PDLVT


MACRO NR2D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END NR2D3BWP240H8P57PDLVT


MACRO INR2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END INR2D1BWP240H8P57PDLVT


MACRO ND2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END ND2D2BWP240H8P57PDLVT


MACRO AO211D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AO211D1BWP240H8P57PDSVT


MACRO IOA21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END IOA21D2BWP240H8P57PDLVT


MACRO IOA21D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END IOA21D4BWP240H8P57PDLVT


MACRO IOA21D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END IOA21D1BWP240H8P57PDLVT


MACRO AO21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AO21D2BWP240H8P57PDSVT


MACRO IOAI21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOAI21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END IOAI21D1BWP240H8P57PDSVT


MACRO OR2D8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D8BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END OR2D8BWP240H8P57PDLVT


MACRO NR4D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END NR4D2BWP240H8P57PDLVT


MACRO AOI32D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AOI32D1BWP240H8P57PDSVT


MACRO OAI211D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OAI211D1BWP240H8P57PDLVT


MACRO BUFFD10BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD10BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END BUFFD10BWP240H8P57PDSVT


MACRO SDFRPQOPTBCD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBCD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END O1

END SDFRPQOPTBCD2BWP240H8P57PDSVT


MACRO SDFRPQOPTBCD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBCD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END O1

END SDFRPQOPTBCD1BWP240H8P57PDSVT


MACRO SDFRPQOPTBCD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBCD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END O1

END SDFRPQOPTBCD1BWP240H8P57PDLVT


MACRO SDFRPQOPTBBD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBBD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.969 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END O1

END SDFRPQOPTBBD1BWP240H8P57PDLVT


MACRO INR3D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END INR3D1BWP240H8P57PDLVT


MACRO OR3D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OR3D1BWP240H8P57PDLVT


MACRO OR2D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OR2D3BWP240H8P57PDSVT


MACRO OR2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OR2D2BWP240H8P57PDSVT


MACRO OAI222D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END OAI222D1BWP240H8P57PDSVT


MACRO OAI21D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END OAI21D1BWP240H8P57PDLVT


MACRO OAI211OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OAI211OPTPAD1BWP240H8P57PDSVT


MACRO IND3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END IND3D1BWP240H8P57PDSVT


MACRO MUX2D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END MUX2D1BWP240H8P57PDSVT


MACRO IOAI21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOAI21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END IOAI21D2BWP240H8P57PDLVT


MACRO NR2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END NR2D2BWP240H8P57PDLVT


MACRO NR4D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END NR4D1BWP240H8P57PDLVT


MACRO AOI21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AOI21D2BWP240H8P57PDSVT


MACRO ND2OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END ND2OPTPAD1BWP240H8P57PDSVT


MACRO NR2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END NR2D2BWP240H8P57PDSVT


MACRO INVSKFD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVSKFD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END INVSKFD4BWP240H8P57PDSVT


MACRO AOI21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AOI21D2BWP240H8P57PDLVT


MACRO OAI21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OAI21D2BWP240H8P57PDSVT


MACRO ND2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END ND2D1BWP240H8P57PDLVT


MACRO NR2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END NR2D1BWP240H8P57PDLVT


MACRO OR2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OR2D2BWP240H8P57PDLVT


MACRO AIOI21D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AIOI21D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AIOI21D1BWP240H8P57PDLVT


MACRO IOA21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END IOA21D2BWP240H8P57PDSVT


MACRO AOI211D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOI211D1BWP240H8P57PDLVT


MACRO XOR2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END XOR2D4BWP240H8P57PDSVT


MACRO OAOI211D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END OAOI211D2BWP240H8P57PDLVT


MACRO SDFSRPQOPTBCD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQOPTBCD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.969 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END O1

END SDFSRPQOPTBCD2BWP240H8P57PDSVT


MACRO OR3D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OR3D2BWP240H8P57PDSVT


MACRO INVPADD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVPADD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END INVPADD1BWP240H8P57PDSVT


MACRO INR4D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR4D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END INR4D1BWP240H8P57PDSVT


MACRO OR2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END OR2D1BWP240H8P57PDLVT


MACRO XOR2D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END XOR2D3BWP240H8P57PDSVT


MACRO ND2OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END ND2OPTPAD1BWP240H8P57PDLVT


MACRO SDFSRPQD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.969 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END O1

END SDFSRPQD1BWP240H8P57PDSVT


MACRO AN4D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN4D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AN4D1BWP240H8P57PDLVT


MACRO ND2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END ND2D2BWP240H8P57PDSVT


MACRO IOA21D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END IOA21D4BWP240H8P57PDSVT


MACRO OAI22D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OAI22D1BWP240H8P57PDLVT


MACRO OAI21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OAI21D2BWP240H8P57PDLVT


MACRO AO22D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AO22D1BWP240H8P57PDLVT


MACRO OAI211D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END OAI211D2BWP240H8P57PDSVT


MACRO ND2D12BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D12BWP240H8P57PDSVT 0 0 ;
  SIZE 1.482 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END O1

END ND2D12BWP240H8P57PDSVT


MACRO OA211D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OA211D1BWP240H8P57PDSVT


MACRO NR2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END NR2D4BWP240H8P57PDSVT


MACRO IIND3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IIND3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END IIND3D1BWP240H8P57PDSVT


MACRO IAO21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAO21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END IAO21D2BWP240H8P57PDSVT


MACRO AO22D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END AO22D2BWP240H8P57PDSVT


MACRO OIAI21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OIAI21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END OIAI21D2BWP240H8P57PDSVT


MACRO NR3D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END NR3D2BWP240H8P57PDSVT


MACRO IAO21D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAO21D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END IAO21D1BWP240H8P57PDLVT


MACRO NR2D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END NR2D3BWP240H8P57PDSVT


MACRO AO211D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AO211D1BWP240H8P57PDLVT


MACRO ND2D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END ND2D4BWP240H8P57PDLVT


MACRO IOA21D6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D6BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END IOA21D6BWP240H8P57PDLVT


MACRO INVD6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END INVD6BWP240H8P57PDLVT


MACRO AOI211OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AOI211OPTPAD1BWP240H8P57PDLVT


MACRO INVD5BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD5BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END INVD5BWP240H8P57PDSVT


MACRO AOI21D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END AOI21D1BWP240H8P57PDLVT


MACRO ND3OPTPAD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3OPTPAD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END ND3OPTPAD2BWP240H8P57PDLVT


MACRO IAO21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAO21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END IAO21D2BWP240H8P57PDLVT


MACRO IINR3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IINR3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END IINR3D1BWP240H8P57PDSVT


MACRO ND4D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END ND4D2BWP240H8P57PDLVT


MACRO AO22D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END AO22D2BWP240H8P57PDLVT


MACRO AN2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END AN2D1BWP240H8P57PDLVT


MACRO INR3OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END INR3OPTPAD1BWP240H8P57PDSVT


MACRO NR2OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END NR2OPTPAD1BWP240H8P57PDLVT


MACRO INVD8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD8BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END INVD8BWP240H8P57PDLVT


MACRO INVD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END INVD4BWP240H8P57PDLVT


MACRO AO22D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END AO22D4BWP240H8P57PDLVT


MACRO IND2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END IND2D1BWP240H8P57PDLVT


MACRO IND2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END IND2D2BWP240H8P57PDSVT


MACRO BUFFSKFD3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END BUFFSKFD3BWP240H8P57PDLVT


MACRO ND2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END ND2D4BWP240H8P57PDSVT


MACRO INVD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.171 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0855 0.12 0.0855 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0855 0.12 0.0855 0.12 ;
    END
  END O1

END INVD1BWP240H8P57PDLVT


MACRO AN3D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN3D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AN3D1BWP240H8P57PDSVT


MACRO AOI21D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END AOI21D4BWP240H8P57PDLVT


MACRO AN2D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AN2D2BWP240H8P57PDSVT


MACRO AOAI211D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END AOAI211D4BWP240H8P57PDLVT


MACRO NR3D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END NR3D2BWP240H8P57PDLVT


MACRO INR3D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END INR3D3BWP240H8P57PDSVT


MACRO INVD3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END INVD3BWP240H8P57PDLVT


MACRO MUX2ND1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2ND1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END MUX2ND1BWP240H8P57PDSVT


MACRO SDFSRPQOPTBBD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQOPTBBD1BWP240H8P57PDSVT 0 0 ;
  SIZE 1.14 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END O1

END SDFSRPQOPTBBD1BWP240H8P57PDSVT


MACRO SDFSRPQOPTBBD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQOPTBBD2BWP240H8P57PDSVT 0 0 ;
  SIZE 1.14 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END O1

END SDFSRPQOPTBBD2BWP240H8P57PDSVT


MACRO SDFSRPQD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.969 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.24 0.4845 0.24 ;
    END
  END O1

END SDFSRPQD1BWP240H8P57PDLVT


MACRO SDFSRPQOPTBBD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQOPTBBD2BWP240H8P57PDLVT 0 0 ;
  SIZE 1.14 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.24 0.57 0.24 ;
    END
  END O1

END SDFSRPQOPTBBD2BWP240H8P57PDLVT


MACRO SDFSRPQOPTBCD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQOPTBCD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.969 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END O1

END SDFSRPQOPTBCD1BWP240H8P57PDLVT


MACRO SDFSRPQOPTBCD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFSRPQOPTBCD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.969 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.36 0.4845 0.36 ;
    END
  END O1

END SDFSRPQOPTBCD2BWP240H8P57PDLVT


MACRO INVD8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD8BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END INVD8BWP240H8P57PDSVT


MACRO AN4D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN4D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AN4D1BWP240H8P57PDSVT


MACRO BUFFSKFD6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END BUFFSKFD6BWP240H8P57PDLVT


MACRO BUFFD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END BUFFD1BWP240H8P57PDLVT


MACRO NR3OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END NR3OPTPAD1BWP240H8P57PDLVT


MACRO AOAI211D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END AOAI211D2BWP240H8P57PDLVT


MACRO ND3D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END ND3D3BWP240H8P57PDLVT


MACRO OA21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OA21D2BWP240H8P57PDLVT


MACRO BUFFD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END BUFFD2BWP240H8P57PDLVT


MACRO MAOI222D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAOI222D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END O1

END MAOI222D2BWP240H8P57PDLVT


MACRO ND2D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND2D3BWP240H8P57PDLVT


MACRO ND3D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END ND3D1BWP240H8P57PDLVT


MACRO NR3OPTPAD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3OPTPAD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END NR3OPTPAD2BWP240H8P57PDLVT


MACRO NR2D6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END NR2D6BWP240H8P57PDSVT


MACRO NR2OPTPAD6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2OPTPAD6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.969 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END O1

END NR2OPTPAD6BWP240H8P57PDSVT


MACRO BUFFD16BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD16BWP240H8P57PDSVT 0 0 ;
  SIZE 0.741 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END O1

END BUFFD16BWP240H8P57PDSVT


MACRO AO21D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.741 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END O1

END AO21D4BWP240H8P57PDSVT


MACRO IOA21D8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D8BWP240H8P57PDLVT 0 0 ;
  SIZE 1.368 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END O1

END IOA21D8BWP240H8P57PDLVT


MACRO ND2SKFD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2SKFD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END ND2SKFD2BWP240H8P57PDLVT


MACRO ND3D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND3D2BWP240H8P57PDLVT


MACRO NR4D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END O1

END NR4D3BWP240H8P57PDSVT


MACRO NR4D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END NR4D2BWP240H8P57PDSVT


MACRO AO22D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END AO22D4BWP240H8P57PDSVT


MACRO ND3OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END ND3OPTPAD1BWP240H8P57PDLVT


MACRO BUFFSKFD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END BUFFSKFD2BWP240H8P57PDLVT


MACRO ND2SKFD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2SKFD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END ND2SKFD4BWP240H8P57PDLVT


MACRO NR4D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END O1

END NR4D3BWP240H8P57PDLVT


MACRO IND4D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND4D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END IND4D1BWP240H8P57PDSVT


MACRO BUFFD14BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD14BWP240H8P57PDSVT 0 0 ;
  SIZE 1.197 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.12 0.5985 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5985 0.12 0.5985 0.12 ;
    END
  END O1

END BUFFD14BWP240H8P57PDSVT


MACRO MUX2D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.741 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END O1

END MUX2D3BWP240H8P57PDSVT


MACRO BUFFD12BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD12BWP240H8P57PDSVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END BUFFD12BWP240H8P57PDSVT


MACRO BUFFD12BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD12BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END BUFFD12BWP240H8P57PDLVT


MACRO AN2D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AN2D3BWP240H8P57PDSVT


MACRO AN2D8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D8BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END AN2D8BWP240H8P57PDSVT


MACRO BUFFD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END BUFFD4BWP240H8P57PDLVT


MACRO BUFFD3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END BUFFD3BWP240H8P57PDLVT


MACRO NR3OPTPAD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3OPTPAD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END NR3OPTPAD4BWP240H8P57PDLVT


MACRO NR2D6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END NR2D6BWP240H8P57PDLVT


MACRO BUFFD10BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD10BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END BUFFD10BWP240H8P57PDLVT


MACRO BUFFSKFD5BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD5BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END BUFFSKFD5BWP240H8P57PDLVT


MACRO AN2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AN2D2BWP240H8P57PDLVT


MACRO IAOI21D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAOI21D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.969 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END O1

END IAOI21D4BWP240H8P57PDLVT


MACRO IAOI21D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAOI21D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.969 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END O1

END IAOI21D4BWP240H8P57PDSVT


MACRO AOI21OPTPAD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21OPTPAD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END AOI21OPTPAD2BWP240H8P57PDLVT


MACRO AOI21D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END AOI21D3BWP240H8P57PDLVT


MACRO AOI21SKFD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21SKFD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END AOI21SKFD4BWP240H8P57PDLVT


MACRO AOI21D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END AOI21D4BWP240H8P57PDSVT


MACRO AOI21OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END AOI21OPTPAD2BWP240H8P57PDSVT


MACRO AOI21D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END AOI21D3BWP240H8P57PDSVT


MACRO IAOI21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAOI21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END IAOI21D2BWP240H8P57PDSVT


MACRO AOI21SKFD6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21SKFD6BWP240H8P57PDSVT 0 0 ;
  SIZE 1.14 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END O1

END AOI21SKFD6BWP240H8P57PDSVT


MACRO ND2SKFD3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2SKFD3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND2SKFD3BWP240H8P57PDLVT


MACRO ND2D6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END ND2D6BWP240H8P57PDSVT


MACRO ND3OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END ND3OPTPAD1BWP240H8P57PDSVT


MACRO FA1D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA1D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END FA1D1BWP240H8P57PDSVT


MACRO IAO22D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAO22D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END IAO22D1BWP240H8P57PDSVT


MACRO INR3OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END INR3OPTPAD2BWP240H8P57PDSVT


MACRO AN3D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN3D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AN3D2BWP240H8P57PDLVT


MACRO INR3D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END INR3D3BWP240H8P57PDLVT


MACRO OR2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END OR2D4BWP240H8P57PDSVT


MACRO IND2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END IND2D2BWP240H8P57PDLVT


MACRO AOAI211D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END AOAI211D1BWP240H8P57PDLVT


MACRO INR2D6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END INR2D6BWP240H8P57PDSVT


MACRO AN4D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN4D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AN4D2BWP240H8P57PDSVT


MACRO ND2D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND2D3BWP240H8P57PDSVT


MACRO OAOI211D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OAOI211D1BWP240H8P57PDLVT


MACRO BUFFD6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END BUFFD6BWP240H8P57PDSVT


MACRO AO211D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END AO211D2BWP240H8P57PDSVT


MACRO OAI211D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END OAI211D2BWP240H8P57PDLVT


MACRO OR4D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OR4D2BWP240H8P57PDLVT


MACRO OAI221D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END OAI221D1BWP240H8P57PDSVT


MACRO NR3D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END NR3D1BWP240H8P57PDLVT


MACRO AN4D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN4D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AN4D2BWP240H8P57PDLVT


MACRO OAI31D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END OAI31D1BWP240H8P57PDLVT


MACRO AIOI21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AIOI21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AIOI21D1BWP240H8P57PDSVT


MACRO OAI211OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END O1

END OAI211OPTPAD2BWP240H8P57PDSVT


MACRO IOA22D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA22D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END IOA22D1BWP240H8P57PDSVT


MACRO IND2D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END IND2D3BWP240H8P57PDLVT


MACRO OIAI21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OIAI21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OIAI21D1BWP240H8P57PDSVT


MACRO ND3D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END ND3D3BWP240H8P57PDSVT


MACRO OAI211SKFD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211SKFD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END OAI211SKFD2BWP240H8P57PDLVT


MACRO AOI222D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END AOI222D1BWP240H8P57PDSVT


MACRO OR2D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END OR2D4BWP240H8P57PDLVT


MACRO BUFFSKFD8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD8BWP240H8P57PDSVT 0 0 ;
  SIZE 0.741 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END O1

END BUFFSKFD8BWP240H8P57PDSVT


MACRO ND3SKFD3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3SKFD3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END ND3SKFD3BWP240H8P57PDLVT


MACRO AOI22OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END AOI22OPTPAD1BWP240H8P57PDLVT


MACRO AOI22D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END AOI22D2BWP240H8P57PDLVT


MACRO BUFFSKFD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END BUFFSKFD4BWP240H8P57PDSVT


MACRO AIOI21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AIOI21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END AIOI21D2BWP240H8P57PDLVT


MACRO IND2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END IND2D4BWP240H8P57PDSVT


MACRO INVD6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END INVD6BWP240H8P57PDSVT


MACRO OA22D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OA22D1BWP240H8P57PDLVT


MACRO OA22D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OA22D1BWP240H8P57PDSVT


MACRO ND3D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND3D2BWP240H8P57PDSVT


MACRO INR3OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END INR3OPTPAD1BWP240H8P57PDLVT


MACRO AOI211D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END AOI211D2BWP240H8P57PDLVT


MACRO AN2D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END AN2D4BWP240H8P57PDLVT


MACRO BUFFSKFD5BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD5BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END BUFFSKFD5BWP240H8P57PDSVT


MACRO IND3D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND3D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END IND3D1BWP240H8P57PDLVT


MACRO BUFFSKFD3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END BUFFSKFD3BWP240H8P57PDSVT


MACRO IND2OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END IND2OPTPAD2BWP240H8P57PDSVT


MACRO INVSKFD3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVSKFD3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.285 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.12 0.1425 0.12 ;
    END
  END O1

END INVSKFD3BWP240H8P57PDSVT


MACRO OAI22D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END OAI22D2BWP240H8P57PDSVT


MACRO ND3OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END ND3OPTPAD2BWP240H8P57PDSVT


MACRO IAOI21D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAOI21D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END IAOI21D2BWP240H8P57PDLVT


MACRO AOI22OPTPAD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22OPTPAD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END O1

END AOI22OPTPAD2BWP240H8P57PDLVT


MACRO ND4SKFD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4SKFD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END ND4SKFD4BWP240H8P57PDSVT


MACRO AN3D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN3D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AN3D1BWP240H8P57PDLVT


MACRO ND2D6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END ND2D6BWP240H8P57PDLVT


MACRO INR3D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END INR3D2BWP240H8P57PDLVT


MACRO INR3OPTPAD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3OPTPAD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END INR3OPTPAD2BWP240H8P57PDLVT


MACRO NR3OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END NR3OPTPAD1BWP240H8P57PDSVT


MACRO ND2SKFD6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2SKFD6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END ND2SKFD6BWP240H8P57PDLVT


MACRO BUFFD6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END BUFFD6BWP240H8P57PDLVT


MACRO BUFFSKFD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END BUFFSKFD4BWP240H8P57PDLVT


MACRO BUFFSKFD8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD8BWP240H8P57PDLVT 0 0 ;
  SIZE 0.741 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.12 0.3705 0.12 ;
    END
  END O1

END BUFFSKFD8BWP240H8P57PDLVT


MACRO OAI21OPTPAD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21OPTPAD4BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END OAI21OPTPAD4BWP240H8P57PDLVT


MACRO INVD5BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVD5BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END INVD5BWP240H8P57PDLVT


MACRO AO21D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AO21D1BWP240H8P57PDSVT


MACRO INR3D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3D4BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END INR3D4BWP240H8P57PDLVT


MACRO NR3OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END NR3OPTPAD2BWP240H8P57PDSVT


MACRO NR2D10BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D10BWP240H8P57PDSVT 0 0 ;
  SIZE 1.254 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END O1

END NR2D10BWP240H8P57PDSVT


MACRO NR2D10BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D10BWP240H8P57PDLVT 0 0 ;
  SIZE 1.254 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END O1

END NR2D10BWP240H8P57PDLVT


MACRO NR2D8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D8BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END NR2D8BWP240H8P57PDLVT


MACRO AOAI211D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END AOAI211D2BWP240H8P57PDSVT


MACRO IND2D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END IND2D4BWP240H8P57PDLVT


MACRO INR2D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END INR2D3BWP240H8P57PDLVT


MACRO XNR2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNR2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END XNR2D4BWP240H8P57PDSVT


MACRO OAOI211D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END OAOI211D4BWP240H8P57PDSVT


MACRO IAOI21D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAOI21D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END IAOI21D1BWP240H8P57PDLVT


MACRO OR4D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OR4D2BWP240H8P57PDSVT


MACRO FCISD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FCISD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END FCISD2BWP240H8P57PDLVT


MACRO INR2OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END INR2OPTPAD1BWP240H8P57PDSVT


MACRO NR2OPTPAD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2OPTPAD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END NR2OPTPAD4BWP240H8P57PDSVT


MACRO INVSKFD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVSKFD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.228 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.12 0.114 0.12 ;
    END
  END O1

END INVSKFD2BWP240H8P57PDSVT


MACRO ND4SKFD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4SKFD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END ND4SKFD2BWP240H8P57PDLVT


MACRO ND3SKFD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3SKFD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND3SKFD2BWP240H8P57PDSVT


MACRO ND3SKFD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3SKFD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END ND3SKFD2BWP240H8P57PDLVT


MACRO INR3OPTPAD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR3OPTPAD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END INR3OPTPAD4BWP240H8P57PDSVT


MACRO SDFRPQOPTBBD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBBD2BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.24 0.513 0.24 ;
    END
  END O1

END SDFRPQOPTBBD2BWP240H8P57PDLVT


MACRO INR2D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END INR2D2BWP240H8P57PDLVT


MACRO IND4D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND4D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END IND4D1BWP240H8P57PDLVT


MACRO OAI211OPTPAD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211OPTPAD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END O1

END OAI211OPTPAD2BWP240H8P57PDLVT


MACRO OAI31D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END OAI31D2BWP240H8P57PDLVT


MACRO AO211D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END AO211D4BWP240H8P57PDLVT


MACRO AOI311D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI311D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AOI311D1BWP240H8P57PDSVT


MACRO OAI311D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI311D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END OAI311D1BWP240H8P57PDSVT


MACRO OAI21D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END OAI21D4BWP240H8P57PDLVT


MACRO INR2OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END INR2OPTPAD2BWP240H8P57PDSVT


MACRO AN3D8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN3D8BWP240H8P57PDSVT 0 0 ;
  SIZE 1.083 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.12 0.5415 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.12 0.5415 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.12 0.5415 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5415 0.12 0.5415 0.12 ;
    END
  END O1

END AN3D8BWP240H8P57PDSVT


MACRO SDFRPQOPTBCD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFRPQOPTBCD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.72 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.36 0.456 0.36 ;
    END
  END O1

END SDFRPQOPTBCD2BWP240H8P57PDLVT


MACRO AOI211OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END O1

END AOI211OPTPAD2BWP240H8P57PDSVT


MACRO FA1D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA1D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END FA1D1BWP240H8P57PDLVT


MACRO XOR2D6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2D6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.741 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END O1

END XOR2D6BWP240H8P57PDLVT


MACRO FCISND1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FCISND1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END FCISND1BWP240H8P57PDSVT


MACRO FCICOD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FCICOD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END FCICOD2BWP240H8P57PDSVT


MACRO ND2SKFD10BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2SKFD10BWP240H8P57PDLVT 0 0 ;
  SIZE 1.254 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.12 0.627 0.12 ;
    END
  END O1

END ND2SKFD10BWP240H8P57PDLVT


MACRO OAI21D8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D8BWP240H8P57PDLVT 0 0 ;
  SIZE 1.482 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END O1

END OAI21D8BWP240H8P57PDLVT


MACRO OAI21D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END OAI21D3BWP240H8P57PDLVT


MACRO ND2D8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D8BWP240H8P57PDSVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END ND2D8BWP240H8P57PDSVT


MACRO FA1OPTCD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA1OPTCD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.24 0.342 0.24 ;
    END
  END O1

END FA1OPTCD1BWP240H8P57PDSVT


MACRO FA1OPTCD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA1OPTCD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.741 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END O1

END FA1OPTCD2BWP240H8P57PDSVT


MACRO HA1D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA1D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END HA1D1BWP240H8P57PDSVT


MACRO FCISD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FCISD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END FCISD2BWP240H8P57PDSVT


MACRO FA1OPTCD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA1OPTCD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.741 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END O1

END FA1OPTCD2BWP240H8P57PDLVT


MACRO FCICOD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FCICOD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END FCICOD1BWP240H8P57PDLVT


MACRO HA1D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA1D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END HA1D2BWP240H8P57PDSVT


MACRO AOI33D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END AOI33D1BWP240H8P57PDSVT


MACRO OR4D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OR4D1BWP240H8P57PDSVT


MACRO AN2D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END AN2D4BWP240H8P57PDSVT


MACRO AN2D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END AN2D3BWP240H8P57PDLVT


MACRO AN2D6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AN2D6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END AN2D6BWP240H8P57PDLVT


MACRO INR2D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END INR2D4BWP240H8P57PDLVT


MACRO INR2D6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INR2D6BWP240H8P57PDLVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END INR2D6BWP240H8P57PDLVT


MACRO AOI222D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.855 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END O1

END AOI222D4BWP240H8P57PDSVT


MACRO IND3D6BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND3D6BWP240H8P57PDLVT 0 0 ;
  SIZE 1.425 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7125 0.12 0.7125 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7125 0.12 0.7125 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7125 0.12 0.7125 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7125 0.12 0.7125 0.12 ;
    END
  END O1

END IND3D6BWP240H8P57PDLVT


MACRO IOA21D8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D8BWP240H8P57PDSVT 0 0 ;
  SIZE 1.368 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.12 0.684 0.12 ;
    END
  END O1

END IOA21D8BWP240H8P57PDSVT


MACRO AOI222D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.24 0.2565 0.24 ;
    END
  END O1

END AOI222D2BWP240H8P57PDLVT


MACRO IND2OPTPAD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND2OPTPAD4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.12 0.456 0.12 ;
    END
  END O1

END IND2OPTPAD4BWP240H8P57PDSVT


MACRO AOI22D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END AOI22D2BWP240H8P57PDSVT


MACRO AOI211D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END AOI211D2BWP240H8P57PDSVT


MACRO AOI222D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.855 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4275 0.24 0.4275 0.24 ;
    END
  END O1

END AOI222D4BWP240H8P57PDLVT


MACRO AOI221D1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221D1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END AOI221D1BWP240H8P57PDSVT


MACRO AOI222D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END AOI222D1BWP240H8P57PDLVT


MACRO ND4SKFD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND4SKFD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.342 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.24 0.171 0.24 ;
    END
  END O1

END ND4SKFD2BWP240H8P57PDSVT


MACRO ND2D8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND2D8BWP240H8P57PDLVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END ND2D8BWP240H8P57PDLVT


MACRO OR4D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.24 0.228 0.24 ;
    END
  END O1

END OR4D4BWP240H8P57PDLVT


MACRO IOAI21D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOAI21D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END IOAI21D1BWP240H8P57PDLVT


MACRO INVSKFD6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVSKFD6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END INVSKFD6BWP240H8P57PDSVT


MACRO ND3D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END ND3D4BWP240H8P57PDLVT


MACRO AOI22OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END AOI22OPTPAD1BWP240H8P57PDSVT


MACRO IOA22D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA22D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END IOA22D1BWP240H8P57PDLVT


MACRO ND3SKFD3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3SKFD3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END ND3SKFD3BWP240H8P57PDSVT


MACRO AOI211OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END AOI211OPTPAD1BWP240H8P57PDSVT


MACRO INVSKFD12BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVSKFD12BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END INVSKFD12BWP240H8P57PDLVT


MACRO BUFFSKFD6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFSKFD6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END BUFFSKFD6BWP240H8P57PDSVT


MACRO ND3SKFD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ND3SKFD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END ND3SKFD4BWP240H8P57PDLVT


MACRO IAO21D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IAO21D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END IAO21D4BWP240H8P57PDLVT


MACRO OAI221D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.399 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.24 0.1995 0.24 ;
    END
  END O1

END OAI221D2BWP240H8P57PDLVT


MACRO OAI221D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I5

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END OAI221D1BWP240H8P57PDLVT


MACRO OA21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OA21D2BWP240H8P57PDSVT


MACRO AOI21D6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D6BWP240H8P57PDSVT 0 0 ;
  SIZE 1.14 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END O1

END AOI21D6BWP240H8P57PDSVT


MACRO AOI21OPTPAD4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21OPTPAD4BWP240H8P57PDSVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END AOI21OPTPAD4BWP240H8P57PDSVT


MACRO IOA22D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA22D4BWP240H8P57PDSVT 0 0 ;
  SIZE 1.14 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.57 0.12 0.57 0.12 ;
    END
  END O1

END IOA22D4BWP240H8P57PDSVT


MACRO OAI31D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END OAI31D4BWP240H8P57PDSVT


MACRO OAI21D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END OAI21D3BWP240H8P57PDSVT


MACRO OAI21OPTPAD2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21OPTPAD2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END OAI21OPTPAD2BWP240H8P57PDLVT


MACRO NR4D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END NR4D4BWP240H8P57PDLVT


MACRO NR3D3BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3D3BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END NR3D3BWP240H8P57PDLVT


MACRO BUFFD16BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFFD16BWP240H8P57PDLVT 0 0 ;
  SIZE 0.741 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3705 0.24 0.3705 0.24 ;
    END
  END O1

END BUFFD16BWP240H8P57PDLVT


MACRO NR4D6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D6BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.24 0.399 0.24 ;
    END
  END O1

END NR4D6BWP240H8P57PDSVT


MACRO NR4D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR4D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END NR4D4BWP240H8P57PDSVT


MACRO INVSKFD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVSKFD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.342 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.12 0.171 0.12 ;
    END
  END O1

END INVSKFD4BWP240H8P57PDLVT


MACRO OAI21D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END OAI21D4BWP240H8P57PDSVT


MACRO IOA21D6BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOA21D6BWP240H8P57PDSVT 0 0 ;
  SIZE 1.026 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.12 0.513 0.12 ;
    END
  END O1

END IOA21D6BWP240H8P57PDSVT


MACRO OAI21OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OAI21OPTPAD1BWP240H8P57PDSVT


MACRO IND3D3BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND3D3BWP240H8P57PDSVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END IND3D3BWP240H8P57PDSVT


MACRO INVSKFD5BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVSKFD5BWP240H8P57PDSVT 0 0 ;
  SIZE 0.399 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END I1

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1995 0.12 0.1995 0.12 ;
    END
  END O1

END INVSKFD5BWP240H8P57PDSVT


MACRO OAI21OPTPAD2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21OPTPAD2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END OAI21OPTPAD2BWP240H8P57PDSVT


MACRO OA211D2BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211D2BWP240H8P57PDLVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END OA211D2BWP240H8P57PDLVT


MACRO OA211D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OA211D1BWP240H8P57PDLVT


MACRO OAI211OPTPAD1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211OPTPAD1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.456 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.12 0.228 0.12 ;
    END
  END O1

END OAI211OPTPAD1BWP240H8P57PDLVT


MACRO OAI222D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I4

  PIN I5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I5

  PIN I6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I6

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END OAI222D1BWP240H8P57PDLVT


MACRO AOI21D8BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21D8BWP240H8P57PDLVT 0 0 ;
  SIZE 1.482 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END O1

END AOI21D8BWP240H8P57PDLVT


MACRO OAI211D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN I4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I4

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END OAI211D4BWP240H8P57PDLVT


MACRO NR3D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.798 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 0.12 0.399 0.12 ;
    END
  END O1

END NR3D4BWP240H8P57PDSVT


MACRO IND3OPTPAD1BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IND3OPTPAD1BWP240H8P57PDSVT 0 0 ;
  SIZE 0.513 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2565 0.12 0.2565 0.12 ;
    END
  END O1

END IND3OPTPAD1BWP240H8P57PDSVT


MACRO MUX2D1BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2D1BWP240H8P57PDLVT 0 0 ;
  SIZE 0.627 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3135 0.12 0.3135 0.12 ;
    END
  END O1

END MUX2D1BWP240H8P57PDLVT


MACRO NR2OPTPAD4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2OPTPAD4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.684 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.12 0.342 0.12 ;
    END
  END O1

END NR2OPTPAD4BWP240H8P57PDLVT


MACRO IOAI21D2BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOAI21D2BWP240H8P57PDSVT 0 0 ;
  SIZE 0.57 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.12 0.285 0.12 ;
    END
  END O1

END IOAI21D2BWP240H8P57PDSVT


MACRO IOAI21D4BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IOAI21D4BWP240H8P57PDSVT 0 0 ;
  SIZE 0.969 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.4845 0.12 0.4845 0.12 ;
    END
  END O1

END IOAI21D4BWP240H8P57PDSVT


MACRO NR3OPTPAD8BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR3OPTPAD8BWP240H8P57PDSVT 0 0 ;
  SIZE 0.912 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.24 0.456 0.24 ;
    END
  END O1

END NR3OPTPAD8BWP240H8P57PDSVT


MACRO IIND3D4BWP240H8P57PDLVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN IIND3D4BWP240H8P57PDLVT 0 0 ;
  SIZE 0.57 BY 0.48 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I2

  PIN I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END I3

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.24 0.285 0.24 ;
    END
  END O1

END IIND3D4BWP240H8P57PDLVT


MACRO NR2D12BWP240H8P57PDSVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NR2D12BWP240H8P57PDSVT 0 0 ;
  SIZE 1.482 BY 0.24 ;
  SYMMETRY Y ;
  SITE FAKE_SITE_1H ;

  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I1

  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END I2

  PIN O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.741 0.12 0.741 0.12 ;
    END
  END O1

END NR2D12BWP240H8P57PDSVT


MACRO sacrls0g4l1p256x16m2b1w0c0p1d0l1rm3sdrw00
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sacrls0g4l1p256x16m2b1w0c0p1d0l1rm3sdrw00 0 0 ;
  SIZE 29.355 BY 19.26 ;
  SYMMETRY X Y ;
  PIN ADR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 15.16 0.342 15.16 ;
    END
  END ADR[0]
  PIN ADR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 15.84 0.171 15.84 ;
    END
  END ADR[1]
  PIN ADR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 16.7915 0.399 16.7915 ;
    END
  END ADR[2]
  PIN ADR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 18.52 0.342 18.52 ;
    END
  END ADR[3]
  PIN ADR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 17.48 0.228 17.48 ;
    END
  END ADR[4]
  PIN ADR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 17.52 0.171 17.52 ;
    END
  END ADR[5]
  PIN ADR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 17.96 0.342 17.96 ;
    END
  END ADR[6]
  PIN ADR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2845 18.0 0.2845 18.0 ;
    END
  END ADR[7]
  PIN BC0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 11.191 0.399 11.191 ;
    END
  END BC0
  PIN BC1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 14.72 0.171 14.72 ;
    END
  END BC1
  PIN BC2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 13.64 0.114 13.64 ;
    END
  END BC2
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 18.04 0.228 18.04 ;
    END
  END CLK
  PIN DFTCLKEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 12.92 0.342 12.92 ;
    END
  END DFTCLKEN
  PIN DFTMASK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 13.08 0.114 13.08 ;
    END
  END DFTMASK
  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 11.96 0.114 11.96 ;
    END
  END DS
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 10.2 0.114 10.2 ;
    END
  END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 4.2 0.114 4.2 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 3.64 0.114 3.64 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 3.0 0.114 3.0 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 2.44 0.114 2.44 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 1.8 0.114 1.8 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 1.24 0.114 1.24 ;
    END
  END D[15]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 9.64 0.114 9.64 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 9.0 0.114 9.0 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 8.44 0.114 8.44 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 7.8 0.114 7.8 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 7.24 0.114 7.24 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 6.6 0.114 6.6 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 6.04 0.114 6.04 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 5.4 0.114 5.4 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 4.84 0.114 4.84 ;
    END
  END D[9]
  PIN FISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 14.6 0.342 14.6 ;
    END
  END FISO
  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2845 17.44 0.2845 17.44 ;
    END
  END LS
  PIN ME
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 11.7515 0.399 11.7515 ;
    END
  END ME
  PIN PIPEME
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 13.04 0.171 13.04 ;
    END
  END PIPEME
  PIN RME
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 12.36 0.342 12.36 ;
    END
  END RME
  PIN RM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 12.48 0.171 12.48 ;
    END
  END RM[0]
  PIN RM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2845 12.4 0.2845 12.4 ;
    END
  END RM[1]
  PIN RM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 12.44 0.228 12.44 ;
    END
  END RM[2]
  PIN RM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 11.8 0.342 11.8 ;
    END
  END RM[3]
  PIN RSCEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 14.04 0.342 14.04 ;
    END
  END RSCEN
  PIN RSCIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 14.68 0.228 14.68 ;
    END
  END RSCIN
  PIN RSCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 14.2 0.114 14.2 ;
    END
  END RSCLK
  PIN RSCRST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 14.12 0.228 14.12 ;
    END
  END RSCRST
  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 13.48 0.342 13.48 ;
    END
  END SD
  PIN SE_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 16.44 0.114 16.44 ;
    END
  END SE_IN
  PIN SE_Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 12.8715 0.399 12.8715 ;
    END
  END SE_Q
  PIN SI_CNTR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 13.4315 0.399 13.4315 ;
    END
  END SI_CNTR
  PIN SI_D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2845 11.84 0.2845 11.84 ;
    END
  END SI_D
  PIN SI_Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 11.88 0.228 11.88 ;
    END
  END SI_Q
  PIN TEST1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 18.68 0.114 18.68 ;
    END
  END TEST1
  PIN TEST_RNM
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2845 12.96 0.2845 12.96 ;
    END
  END TEST_RNM
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 18.64 0.171 18.64 ;
    END
  END WE
  PIN QP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 10.12 0.228 10.12 ;
    END
  END QP[0]
  PIN QP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 4.12 0.228 4.12 ;
    END
  END QP[10]
  PIN QP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 3.56 0.228 3.56 ;
    END
  END QP[11]
  PIN QP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 2.92 0.228 2.92 ;
    END
  END QP[12]
  PIN QP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 2.36 0.228 2.36 ;
    END
  END QP[13]
  PIN QP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 1.72 0.228 1.72 ;
    END
  END QP[14]
  PIN QP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 1.16 0.228 1.16 ;
    END
  END QP[15]
  PIN QP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 9.56 0.228 9.56 ;
    END
  END QP[1]
  PIN QP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 8.92 0.228 8.92 ;
    END
  END QP[2]
  PIN QP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 8.36 0.228 8.36 ;
    END
  END QP[3]
  PIN QP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 7.72 0.228 7.72 ;
    END
  END QP[4]
  PIN QP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 7.16 0.228 7.16 ;
    END
  END QP[5]
  PIN QP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 6.52 0.228 6.52 ;
    END
  END QP[6]
  PIN QP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 5.96 0.228 5.96 ;
    END
  END QP[7]
  PIN QP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 5.32 0.228 5.32 ;
    END
  END QP[8]
  PIN QP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 4.76 0.228 4.76 ;
    END
  END QP[9]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 10.16 0.171 10.16 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 4.16 0.171 4.16 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 3.6 0.171 3.6 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 2.96 0.171 2.96 ;
    END
  END Q[12]
  PIN Q[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 2.4 0.171 2.4 ;
    END
  END Q[13]
  PIN Q[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 1.76 0.171 1.76 ;
    END
  END Q[14]
  PIN Q[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 1.2 0.171 1.2 ;
    END
  END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 9.6 0.171 9.6 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 8.96 0.171 8.96 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 8.4 0.171 8.4 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 7.76 0.171 7.76 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 7.2 0.171 7.2 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 6.56 0.171 6.56 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 6.0 0.171 6.0 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 5.36 0.171 5.36 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 4.8 0.171 4.8 ;
    END
  END Q[9]
  PIN ROP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.5 0.171 0.5 ;
    END
  END ROP
  PIN RSCOUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.399 13.992 0.399 13.992 ;
    END
  END RSCOUT
  PIN SO_CNTR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 11.24 0.342 11.24 ;
    END
  END SO_CNTR
  PIN SO_D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.54 0.114 0.54 ;
    END
  END SO_D
  PIN SO_Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.46 0.228 0.46 ;
    END
  END SO_Q
END sacrls0g4l1p256x16m2b1w0c0p1d0l1rm3sdrw00


END LIBRARY