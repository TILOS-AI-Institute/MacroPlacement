VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_256x32
  FOREIGN fakeram130_256x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 293.940 BY 349.520 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 4.370 0.460 4.830 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.130 0.460 7.590 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.890 0.460 10.350 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.650 0.460 13.110 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 15.410 0.460 15.870 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.170 0.460 18.630 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.930 0.460 21.390 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.690 0.460 24.150 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.450 0.460 26.910 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.210 0.460 29.670 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.970 0.460 32.430 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.730 0.460 35.190 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.490 0.460 37.950 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.250 0.460 40.710 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.010 0.460 43.470 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.770 0.460 46.230 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 48.530 0.460 48.990 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 51.290 0.460 51.750 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.050 0.460 54.510 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.810 0.460 57.270 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.570 0.460 60.030 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.330 0.460 62.790 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 65.090 0.460 65.550 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.850 0.460 68.310 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.610 0.460 71.070 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.370 0.460 73.830 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.130 0.460 76.590 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.890 0.460 79.350 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.650 0.460 82.110 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.410 0.460 84.870 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 87.170 0.460 87.630 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.930 0.460 90.390 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.970 0.460 101.430 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.730 0.460 104.190 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.490 0.460 106.950 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 109.250 0.460 109.710 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.010 0.460 112.470 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 114.770 0.460 115.230 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 117.530 0.460 117.990 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.290 0.460 120.750 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.050 0.460 123.510 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 125.810 0.460 126.270 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 128.570 0.460 129.030 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.330 0.460 131.790 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.090 0.460 134.550 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.850 0.460 137.310 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.610 0.460 140.070 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.370 0.460 142.830 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.130 0.460 145.590 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 147.890 0.460 148.350 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.650 0.460 151.110 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.410 0.460 153.870 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.170 0.460 156.630 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.930 0.460 159.390 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.690 0.460 162.150 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.450 0.460 164.910 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.210 0.460 167.670 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.970 0.460 170.430 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 172.730 0.460 173.190 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.490 0.460 175.950 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 178.250 0.460 178.710 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 181.010 0.460 181.470 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 183.770 0.460 184.230 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.530 0.460 186.990 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 197.570 0.460 198.030 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 200.330 0.460 200.790 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 203.090 0.460 203.550 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.850 0.460 206.310 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 208.610 0.460 209.070 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 211.370 0.460 211.830 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 214.130 0.460 214.590 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.890 0.460 217.350 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 219.650 0.460 220.110 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 222.410 0.460 222.870 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 225.170 0.460 225.630 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 227.930 0.460 228.390 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 230.690 0.460 231.150 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 233.450 0.460 233.910 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 236.210 0.460 236.670 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 238.970 0.460 239.430 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 241.730 0.460 242.190 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 244.490 0.460 244.950 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 247.250 0.460 247.710 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 250.010 0.460 250.470 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 252.770 0.460 253.230 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 255.530 0.460 255.990 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 258.290 0.460 258.750 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 261.050 0.460 261.510 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 263.810 0.460 264.270 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 266.570 0.460 267.030 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 269.330 0.460 269.790 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 272.090 0.460 272.550 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 274.850 0.460 275.310 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 277.610 0.460 278.070 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 280.370 0.460 280.830 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 283.130 0.460 283.590 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 294.170 0.460 294.630 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 296.930 0.460 297.390 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 299.690 0.460 300.150 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 302.450 0.460 302.910 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 305.210 0.460 305.670 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 307.970 0.460 308.430 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 310.730 0.460 311.190 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 313.490 0.460 313.950 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 324.530 0.460 324.990 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.290 0.460 327.750 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.050 0.460 330.510 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.680 4.600 5.520 344.920 ;
      RECT 11.040 4.600 12.880 344.920 ;
      RECT 18.400 4.600 20.240 344.920 ;
      RECT 25.760 4.600 27.600 344.920 ;
      RECT 33.120 4.600 34.960 344.920 ;
      RECT 40.480 4.600 42.320 344.920 ;
      RECT 47.840 4.600 49.680 344.920 ;
      RECT 55.200 4.600 57.040 344.920 ;
      RECT 62.560 4.600 64.400 344.920 ;
      RECT 69.920 4.600 71.760 344.920 ;
      RECT 77.280 4.600 79.120 344.920 ;
      RECT 84.640 4.600 86.480 344.920 ;
      RECT 92.000 4.600 93.840 344.920 ;
      RECT 99.360 4.600 101.200 344.920 ;
      RECT 106.720 4.600 108.560 344.920 ;
      RECT 114.080 4.600 115.920 344.920 ;
      RECT 121.440 4.600 123.280 344.920 ;
      RECT 128.800 4.600 130.640 344.920 ;
      RECT 136.160 4.600 138.000 344.920 ;
      RECT 143.520 4.600 145.360 344.920 ;
      RECT 150.880 4.600 152.720 344.920 ;
      RECT 158.240 4.600 160.080 344.920 ;
      RECT 165.600 4.600 167.440 344.920 ;
      RECT 172.960 4.600 174.800 344.920 ;
      RECT 180.320 4.600 182.160 344.920 ;
      RECT 187.680 4.600 189.520 344.920 ;
      RECT 195.040 4.600 196.880 344.920 ;
      RECT 202.400 4.600 204.240 344.920 ;
      RECT 209.760 4.600 211.600 344.920 ;
      RECT 217.120 4.600 218.960 344.920 ;
      RECT 224.480 4.600 226.320 344.920 ;
      RECT 231.840 4.600 233.680 344.920 ;
      RECT 239.200 4.600 241.040 344.920 ;
      RECT 246.560 4.600 248.400 344.920 ;
      RECT 253.920 4.600 255.760 344.920 ;
      RECT 261.280 4.600 263.120 344.920 ;
      RECT 268.640 4.600 270.480 344.920 ;
      RECT 276.000 4.600 277.840 344.920 ;
      RECT 283.360 4.600 285.200 344.920 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 7.360 4.600 9.200 344.920 ;
      RECT 14.720 4.600 16.560 344.920 ;
      RECT 22.080 4.600 23.920 344.920 ;
      RECT 29.440 4.600 31.280 344.920 ;
      RECT 36.800 4.600 38.640 344.920 ;
      RECT 44.160 4.600 46.000 344.920 ;
      RECT 51.520 4.600 53.360 344.920 ;
      RECT 58.880 4.600 60.720 344.920 ;
      RECT 66.240 4.600 68.080 344.920 ;
      RECT 73.600 4.600 75.440 344.920 ;
      RECT 80.960 4.600 82.800 344.920 ;
      RECT 88.320 4.600 90.160 344.920 ;
      RECT 95.680 4.600 97.520 344.920 ;
      RECT 103.040 4.600 104.880 344.920 ;
      RECT 110.400 4.600 112.240 344.920 ;
      RECT 117.760 4.600 119.600 344.920 ;
      RECT 125.120 4.600 126.960 344.920 ;
      RECT 132.480 4.600 134.320 344.920 ;
      RECT 139.840 4.600 141.680 344.920 ;
      RECT 147.200 4.600 149.040 344.920 ;
      RECT 154.560 4.600 156.400 344.920 ;
      RECT 161.920 4.600 163.760 344.920 ;
      RECT 169.280 4.600 171.120 344.920 ;
      RECT 176.640 4.600 178.480 344.920 ;
      RECT 184.000 4.600 185.840 344.920 ;
      RECT 191.360 4.600 193.200 344.920 ;
      RECT 198.720 4.600 200.560 344.920 ;
      RECT 206.080 4.600 207.920 344.920 ;
      RECT 213.440 4.600 215.280 344.920 ;
      RECT 220.800 4.600 222.640 344.920 ;
      RECT 228.160 4.600 230.000 344.920 ;
      RECT 235.520 4.600 237.360 344.920 ;
      RECT 242.880 4.600 244.720 344.920 ;
      RECT 250.240 4.600 252.080 344.920 ;
      RECT 257.600 4.600 259.440 344.920 ;
      RECT 264.960 4.600 266.800 344.920 ;
      RECT 272.320 4.600 274.160 344.920 ;
      RECT 279.680 4.600 281.520 344.920 ;
      RECT 287.040 4.600 288.880 344.920 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 293.940 349.520 ;
    LAYER met2 ;
    RECT 0 0 293.940 349.520 ;
    LAYER met3 ;
    RECT 0.460 0 293.940 349.520 ;
    RECT 0 0.000 0.460 4.370 ;
    RECT 0 4.830 0.460 7.130 ;
    RECT 0 7.590 0.460 9.890 ;
    RECT 0 10.350 0.460 12.650 ;
    RECT 0 13.110 0.460 15.410 ;
    RECT 0 15.870 0.460 18.170 ;
    RECT 0 18.630 0.460 20.930 ;
    RECT 0 21.390 0.460 23.690 ;
    RECT 0 24.150 0.460 26.450 ;
    RECT 0 26.910 0.460 29.210 ;
    RECT 0 29.670 0.460 31.970 ;
    RECT 0 32.430 0.460 34.730 ;
    RECT 0 35.190 0.460 37.490 ;
    RECT 0 37.950 0.460 40.250 ;
    RECT 0 40.710 0.460 43.010 ;
    RECT 0 43.470 0.460 45.770 ;
    RECT 0 46.230 0.460 48.530 ;
    RECT 0 48.990 0.460 51.290 ;
    RECT 0 51.750 0.460 54.050 ;
    RECT 0 54.510 0.460 56.810 ;
    RECT 0 57.270 0.460 59.570 ;
    RECT 0 60.030 0.460 62.330 ;
    RECT 0 62.790 0.460 65.090 ;
    RECT 0 65.550 0.460 67.850 ;
    RECT 0 68.310 0.460 70.610 ;
    RECT 0 71.070 0.460 73.370 ;
    RECT 0 73.830 0.460 76.130 ;
    RECT 0 76.590 0.460 78.890 ;
    RECT 0 79.350 0.460 81.650 ;
    RECT 0 82.110 0.460 84.410 ;
    RECT 0 84.870 0.460 87.170 ;
    RECT 0 87.630 0.460 89.930 ;
    RECT 0 90.390 0.460 100.970 ;
    RECT 0 101.430 0.460 103.730 ;
    RECT 0 104.190 0.460 106.490 ;
    RECT 0 106.950 0.460 109.250 ;
    RECT 0 109.710 0.460 112.010 ;
    RECT 0 112.470 0.460 114.770 ;
    RECT 0 115.230 0.460 117.530 ;
    RECT 0 117.990 0.460 120.290 ;
    RECT 0 120.750 0.460 123.050 ;
    RECT 0 123.510 0.460 125.810 ;
    RECT 0 126.270 0.460 128.570 ;
    RECT 0 129.030 0.460 131.330 ;
    RECT 0 131.790 0.460 134.090 ;
    RECT 0 134.550 0.460 136.850 ;
    RECT 0 137.310 0.460 139.610 ;
    RECT 0 140.070 0.460 142.370 ;
    RECT 0 142.830 0.460 145.130 ;
    RECT 0 145.590 0.460 147.890 ;
    RECT 0 148.350 0.460 150.650 ;
    RECT 0 151.110 0.460 153.410 ;
    RECT 0 153.870 0.460 156.170 ;
    RECT 0 156.630 0.460 158.930 ;
    RECT 0 159.390 0.460 161.690 ;
    RECT 0 162.150 0.460 164.450 ;
    RECT 0 164.910 0.460 167.210 ;
    RECT 0 167.670 0.460 169.970 ;
    RECT 0 170.430 0.460 172.730 ;
    RECT 0 173.190 0.460 175.490 ;
    RECT 0 175.950 0.460 178.250 ;
    RECT 0 178.710 0.460 181.010 ;
    RECT 0 181.470 0.460 183.770 ;
    RECT 0 184.230 0.460 186.530 ;
    RECT 0 186.990 0.460 197.570 ;
    RECT 0 198.030 0.460 200.330 ;
    RECT 0 200.790 0.460 203.090 ;
    RECT 0 203.550 0.460 205.850 ;
    RECT 0 206.310 0.460 208.610 ;
    RECT 0 209.070 0.460 211.370 ;
    RECT 0 211.830 0.460 214.130 ;
    RECT 0 214.590 0.460 216.890 ;
    RECT 0 217.350 0.460 219.650 ;
    RECT 0 220.110 0.460 222.410 ;
    RECT 0 222.870 0.460 225.170 ;
    RECT 0 225.630 0.460 227.930 ;
    RECT 0 228.390 0.460 230.690 ;
    RECT 0 231.150 0.460 233.450 ;
    RECT 0 233.910 0.460 236.210 ;
    RECT 0 236.670 0.460 238.970 ;
    RECT 0 239.430 0.460 241.730 ;
    RECT 0 242.190 0.460 244.490 ;
    RECT 0 244.950 0.460 247.250 ;
    RECT 0 247.710 0.460 250.010 ;
    RECT 0 250.470 0.460 252.770 ;
    RECT 0 253.230 0.460 255.530 ;
    RECT 0 255.990 0.460 258.290 ;
    RECT 0 258.750 0.460 261.050 ;
    RECT 0 261.510 0.460 263.810 ;
    RECT 0 264.270 0.460 266.570 ;
    RECT 0 267.030 0.460 269.330 ;
    RECT 0 269.790 0.460 272.090 ;
    RECT 0 272.550 0.460 274.850 ;
    RECT 0 275.310 0.460 277.610 ;
    RECT 0 278.070 0.460 280.370 ;
    RECT 0 280.830 0.460 283.130 ;
    RECT 0 283.590 0.460 294.170 ;
    RECT 0 294.630 0.460 296.930 ;
    RECT 0 297.390 0.460 299.690 ;
    RECT 0 300.150 0.460 302.450 ;
    RECT 0 302.910 0.460 305.210 ;
    RECT 0 305.670 0.460 307.970 ;
    RECT 0 308.430 0.460 310.730 ;
    RECT 0 311.190 0.460 313.490 ;
    RECT 0 313.950 0.460 324.530 ;
    RECT 0 324.990 0.460 327.290 ;
    RECT 0 327.750 0.460 330.050 ;
    RECT 0 330.510 0.460 349.520 ;
    LAYER met4 ;
    RECT 0 0 293.940 4.600 ;
    RECT 0 344.920 293.940 349.520 ;
    RECT 0.000 4.600 3.680 344.920 ;
    RECT 5.520 4.600 7.360 344.920 ;
    RECT 9.200 4.600 11.040 344.920 ;
    RECT 12.880 4.600 14.720 344.920 ;
    RECT 16.560 4.600 18.400 344.920 ;
    RECT 20.240 4.600 22.080 344.920 ;
    RECT 23.920 4.600 25.760 344.920 ;
    RECT 27.600 4.600 29.440 344.920 ;
    RECT 31.280 4.600 33.120 344.920 ;
    RECT 34.960 4.600 36.800 344.920 ;
    RECT 38.640 4.600 40.480 344.920 ;
    RECT 42.320 4.600 44.160 344.920 ;
    RECT 46.000 4.600 47.840 344.920 ;
    RECT 49.680 4.600 51.520 344.920 ;
    RECT 53.360 4.600 55.200 344.920 ;
    RECT 57.040 4.600 58.880 344.920 ;
    RECT 60.720 4.600 62.560 344.920 ;
    RECT 64.400 4.600 66.240 344.920 ;
    RECT 68.080 4.600 69.920 344.920 ;
    RECT 71.760 4.600 73.600 344.920 ;
    RECT 75.440 4.600 77.280 344.920 ;
    RECT 79.120 4.600 80.960 344.920 ;
    RECT 82.800 4.600 84.640 344.920 ;
    RECT 86.480 4.600 88.320 344.920 ;
    RECT 90.160 4.600 92.000 344.920 ;
    RECT 93.840 4.600 95.680 344.920 ;
    RECT 97.520 4.600 99.360 344.920 ;
    RECT 101.200 4.600 103.040 344.920 ;
    RECT 104.880 4.600 106.720 344.920 ;
    RECT 108.560 4.600 110.400 344.920 ;
    RECT 112.240 4.600 114.080 344.920 ;
    RECT 115.920 4.600 117.760 344.920 ;
    RECT 119.600 4.600 121.440 344.920 ;
    RECT 123.280 4.600 125.120 344.920 ;
    RECT 126.960 4.600 128.800 344.920 ;
    RECT 130.640 4.600 132.480 344.920 ;
    RECT 134.320 4.600 136.160 344.920 ;
    RECT 138.000 4.600 139.840 344.920 ;
    RECT 141.680 4.600 143.520 344.920 ;
    RECT 145.360 4.600 147.200 344.920 ;
    RECT 149.040 4.600 150.880 344.920 ;
    RECT 152.720 4.600 154.560 344.920 ;
    RECT 156.400 4.600 158.240 344.920 ;
    RECT 160.080 4.600 161.920 344.920 ;
    RECT 163.760 4.600 165.600 344.920 ;
    RECT 167.440 4.600 169.280 344.920 ;
    RECT 171.120 4.600 172.960 344.920 ;
    RECT 174.800 4.600 176.640 344.920 ;
    RECT 178.480 4.600 180.320 344.920 ;
    RECT 182.160 4.600 184.000 344.920 ;
    RECT 185.840 4.600 187.680 344.920 ;
    RECT 189.520 4.600 191.360 344.920 ;
    RECT 193.200 4.600 195.040 344.920 ;
    RECT 196.880 4.600 198.720 344.920 ;
    RECT 200.560 4.600 202.400 344.920 ;
    RECT 204.240 4.600 206.080 344.920 ;
    RECT 207.920 4.600 209.760 344.920 ;
    RECT 211.600 4.600 213.440 344.920 ;
    RECT 215.280 4.600 217.120 344.920 ;
    RECT 218.960 4.600 220.800 344.920 ;
    RECT 222.640 4.600 224.480 344.920 ;
    RECT 226.320 4.600 228.160 344.920 ;
    RECT 230.000 4.600 231.840 344.920 ;
    RECT 233.680 4.600 235.520 344.920 ;
    RECT 237.360 4.600 239.200 344.920 ;
    RECT 241.040 4.600 242.880 344.920 ;
    RECT 244.720 4.600 246.560 344.920 ;
    RECT 248.400 4.600 250.240 344.920 ;
    RECT 252.080 4.600 253.920 344.920 ;
    RECT 255.760 4.600 257.600 344.920 ;
    RECT 259.440 4.600 261.280 344.920 ;
    RECT 263.120 4.600 264.960 344.920 ;
    RECT 266.800 4.600 268.640 344.920 ;
    RECT 270.480 4.600 272.320 344.920 ;
    RECT 274.160 4.600 276.000 344.920 ;
    RECT 277.840 4.600 279.680 344.920 ;
    RECT 281.520 4.600 283.360 344.920 ;
    RECT 285.200 4.600 287.040 344.920 ;
    RECT 288.880 4.600 293.940 344.920 ;
    LAYER OVERLAP ;
    RECT 0 0 293.940 349.520 ;
  END
END fakeram130_256x32

END LIBRARY
