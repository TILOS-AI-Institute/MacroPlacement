VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_256x512
  FOREIGN fakeram130_256x512 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 834.440 BY 1052.640 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 4.370 0.460 4.830 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 4.830 0.460 5.290 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.290 0.460 5.750 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.750 0.460 6.210 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.210 0.460 6.670 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.670 0.460 7.130 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.130 0.460 7.590 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.590 0.460 8.050 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.050 0.460 8.510 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.510 0.460 8.970 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.970 0.460 9.430 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.430 0.460 9.890 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.890 0.460 10.350 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.350 0.460 10.810 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.810 0.460 11.270 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 11.270 0.460 11.730 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 11.730 0.460 12.190 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.190 0.460 12.650 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.650 0.460 13.110 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.110 0.460 13.570 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.570 0.460 14.030 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.030 0.460 14.490 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.490 0.460 14.950 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.950 0.460 15.410 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 15.410 0.460 15.870 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 15.870 0.460 16.330 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.330 0.460 16.790 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.790 0.460 17.250 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.250 0.460 17.710 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.710 0.460 18.170 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.170 0.460 18.630 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.630 0.460 19.090 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 19.090 0.460 19.550 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 19.550 0.460 20.010 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.010 0.460 20.470 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.470 0.460 20.930 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.930 0.460 21.390 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.390 0.460 21.850 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.850 0.460 22.310 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.310 0.460 22.770 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.770 0.460 23.230 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.230 0.460 23.690 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.690 0.460 24.150 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.150 0.460 24.610 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.610 0.460 25.070 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.070 0.460 25.530 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.530 0.460 25.990 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.990 0.460 26.450 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.450 0.460 26.910 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.910 0.460 27.370 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.370 0.460 27.830 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.830 0.460 28.290 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.290 0.460 28.750 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.750 0.460 29.210 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.210 0.460 29.670 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.670 0.460 30.130 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 30.130 0.460 30.590 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 30.590 0.460 31.050 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.050 0.460 31.510 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.510 0.460 31.970 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.970 0.460 32.430 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.430 0.460 32.890 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.890 0.460 33.350 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.350 0.460 33.810 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.810 0.460 34.270 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.270 0.460 34.730 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.730 0.460 35.190 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.190 0.460 35.650 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.650 0.460 36.110 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 36.110 0.460 36.570 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 36.570 0.460 37.030 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.030 0.460 37.490 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.490 0.460 37.950 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.950 0.460 38.410 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.410 0.460 38.870 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.870 0.460 39.330 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.330 0.460 39.790 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.790 0.460 40.250 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.250 0.460 40.710 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.710 0.460 41.170 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.170 0.460 41.630 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.630 0.460 42.090 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.090 0.460 42.550 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.550 0.460 43.010 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.010 0.460 43.470 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.470 0.460 43.930 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.930 0.460 44.390 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.390 0.460 44.850 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.850 0.460 45.310 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.310 0.460 45.770 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.770 0.460 46.230 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 46.230 0.460 46.690 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 46.690 0.460 47.150 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.150 0.460 47.610 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.610 0.460 48.070 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 48.070 0.460 48.530 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 48.530 0.460 48.990 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 48.990 0.460 49.450 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 49.450 0.460 49.910 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 49.910 0.460 50.370 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.370 0.460 50.830 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.830 0.460 51.290 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 51.290 0.460 51.750 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 51.750 0.460 52.210 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.210 0.460 52.670 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.670 0.460 53.130 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 53.130 0.460 53.590 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 53.590 0.460 54.050 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.050 0.460 54.510 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.510 0.460 54.970 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.970 0.460 55.430 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.430 0.460 55.890 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.890 0.460 56.350 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.350 0.460 56.810 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.810 0.460 57.270 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 57.270 0.460 57.730 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 57.730 0.460 58.190 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 58.190 0.460 58.650 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 58.650 0.460 59.110 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.110 0.460 59.570 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.570 0.460 60.030 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 60.030 0.460 60.490 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 60.490 0.460 60.950 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 60.950 0.460 61.410 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 61.410 0.460 61.870 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 61.870 0.460 62.330 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.330 0.460 62.790 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.790 0.460 63.250 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.250 0.460 63.710 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.710 0.460 64.170 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.170 0.460 64.630 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.630 0.460 65.090 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 65.090 0.460 65.550 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 65.550 0.460 66.010 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.010 0.460 66.470 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.470 0.460 66.930 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.930 0.460 67.390 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.390 0.460 67.850 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.850 0.460 68.310 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 68.310 0.460 68.770 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 68.770 0.460 69.230 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.230 0.460 69.690 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.690 0.460 70.150 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.150 0.460 70.610 ;
    END
  END w_mask_in[143]
  PIN w_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.610 0.460 71.070 ;
    END
  END w_mask_in[144]
  PIN w_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.070 0.460 71.530 ;
    END
  END w_mask_in[145]
  PIN w_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.530 0.460 71.990 ;
    END
  END w_mask_in[146]
  PIN w_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.990 0.460 72.450 ;
    END
  END w_mask_in[147]
  PIN w_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 72.450 0.460 72.910 ;
    END
  END w_mask_in[148]
  PIN w_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 72.910 0.460 73.370 ;
    END
  END w_mask_in[149]
  PIN w_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.370 0.460 73.830 ;
    END
  END w_mask_in[150]
  PIN w_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.830 0.460 74.290 ;
    END
  END w_mask_in[151]
  PIN w_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.290 0.460 74.750 ;
    END
  END w_mask_in[152]
  PIN w_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.750 0.460 75.210 ;
    END
  END w_mask_in[153]
  PIN w_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 75.210 0.460 75.670 ;
    END
  END w_mask_in[154]
  PIN w_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 75.670 0.460 76.130 ;
    END
  END w_mask_in[155]
  PIN w_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.130 0.460 76.590 ;
    END
  END w_mask_in[156]
  PIN w_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.590 0.460 77.050 ;
    END
  END w_mask_in[157]
  PIN w_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.050 0.460 77.510 ;
    END
  END w_mask_in[158]
  PIN w_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.510 0.460 77.970 ;
    END
  END w_mask_in[159]
  PIN w_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.970 0.460 78.430 ;
    END
  END w_mask_in[160]
  PIN w_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.430 0.460 78.890 ;
    END
  END w_mask_in[161]
  PIN w_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.890 0.460 79.350 ;
    END
  END w_mask_in[162]
  PIN w_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.350 0.460 79.810 ;
    END
  END w_mask_in[163]
  PIN w_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.810 0.460 80.270 ;
    END
  END w_mask_in[164]
  PIN w_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.270 0.460 80.730 ;
    END
  END w_mask_in[165]
  PIN w_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.730 0.460 81.190 ;
    END
  END w_mask_in[166]
  PIN w_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.190 0.460 81.650 ;
    END
  END w_mask_in[167]
  PIN w_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.650 0.460 82.110 ;
    END
  END w_mask_in[168]
  PIN w_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.110 0.460 82.570 ;
    END
  END w_mask_in[169]
  PIN w_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.570 0.460 83.030 ;
    END
  END w_mask_in[170]
  PIN w_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.030 0.460 83.490 ;
    END
  END w_mask_in[171]
  PIN w_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.490 0.460 83.950 ;
    END
  END w_mask_in[172]
  PIN w_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.950 0.460 84.410 ;
    END
  END w_mask_in[173]
  PIN w_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.410 0.460 84.870 ;
    END
  END w_mask_in[174]
  PIN w_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.870 0.460 85.330 ;
    END
  END w_mask_in[175]
  PIN w_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.330 0.460 85.790 ;
    END
  END w_mask_in[176]
  PIN w_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.790 0.460 86.250 ;
    END
  END w_mask_in[177]
  PIN w_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.250 0.460 86.710 ;
    END
  END w_mask_in[178]
  PIN w_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.710 0.460 87.170 ;
    END
  END w_mask_in[179]
  PIN w_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 87.170 0.460 87.630 ;
    END
  END w_mask_in[180]
  PIN w_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 87.630 0.460 88.090 ;
    END
  END w_mask_in[181]
  PIN w_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.090 0.460 88.550 ;
    END
  END w_mask_in[182]
  PIN w_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.550 0.460 89.010 ;
    END
  END w_mask_in[183]
  PIN w_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.010 0.460 89.470 ;
    END
  END w_mask_in[184]
  PIN w_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.470 0.460 89.930 ;
    END
  END w_mask_in[185]
  PIN w_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.930 0.460 90.390 ;
    END
  END w_mask_in[186]
  PIN w_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.390 0.460 90.850 ;
    END
  END w_mask_in[187]
  PIN w_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.850 0.460 91.310 ;
    END
  END w_mask_in[188]
  PIN w_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 91.310 0.460 91.770 ;
    END
  END w_mask_in[189]
  PIN w_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 91.770 0.460 92.230 ;
    END
  END w_mask_in[190]
  PIN w_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.230 0.460 92.690 ;
    END
  END w_mask_in[191]
  PIN w_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.690 0.460 93.150 ;
    END
  END w_mask_in[192]
  PIN w_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.150 0.460 93.610 ;
    END
  END w_mask_in[193]
  PIN w_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.610 0.460 94.070 ;
    END
  END w_mask_in[194]
  PIN w_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.070 0.460 94.530 ;
    END
  END w_mask_in[195]
  PIN w_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.530 0.460 94.990 ;
    END
  END w_mask_in[196]
  PIN w_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.990 0.460 95.450 ;
    END
  END w_mask_in[197]
  PIN w_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.450 0.460 95.910 ;
    END
  END w_mask_in[198]
  PIN w_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.910 0.460 96.370 ;
    END
  END w_mask_in[199]
  PIN w_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.370 0.460 96.830 ;
    END
  END w_mask_in[200]
  PIN w_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.830 0.460 97.290 ;
    END
  END w_mask_in[201]
  PIN w_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.290 0.460 97.750 ;
    END
  END w_mask_in[202]
  PIN w_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.750 0.460 98.210 ;
    END
  END w_mask_in[203]
  PIN w_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 98.210 0.460 98.670 ;
    END
  END w_mask_in[204]
  PIN w_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 98.670 0.460 99.130 ;
    END
  END w_mask_in[205]
  PIN w_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.130 0.460 99.590 ;
    END
  END w_mask_in[206]
  PIN w_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.590 0.460 100.050 ;
    END
  END w_mask_in[207]
  PIN w_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.050 0.460 100.510 ;
    END
  END w_mask_in[208]
  PIN w_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.510 0.460 100.970 ;
    END
  END w_mask_in[209]
  PIN w_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.970 0.460 101.430 ;
    END
  END w_mask_in[210]
  PIN w_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.430 0.460 101.890 ;
    END
  END w_mask_in[211]
  PIN w_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.890 0.460 102.350 ;
    END
  END w_mask_in[212]
  PIN w_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.350 0.460 102.810 ;
    END
  END w_mask_in[213]
  PIN w_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.810 0.460 103.270 ;
    END
  END w_mask_in[214]
  PIN w_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.270 0.460 103.730 ;
    END
  END w_mask_in[215]
  PIN w_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.730 0.460 104.190 ;
    END
  END w_mask_in[216]
  PIN w_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.190 0.460 104.650 ;
    END
  END w_mask_in[217]
  PIN w_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.650 0.460 105.110 ;
    END
  END w_mask_in[218]
  PIN w_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.110 0.460 105.570 ;
    END
  END w_mask_in[219]
  PIN w_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.570 0.460 106.030 ;
    END
  END w_mask_in[220]
  PIN w_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.030 0.460 106.490 ;
    END
  END w_mask_in[221]
  PIN w_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.490 0.460 106.950 ;
    END
  END w_mask_in[222]
  PIN w_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.950 0.460 107.410 ;
    END
  END w_mask_in[223]
  PIN w_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.410 0.460 107.870 ;
    END
  END w_mask_in[224]
  PIN w_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.870 0.460 108.330 ;
    END
  END w_mask_in[225]
  PIN w_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 108.330 0.460 108.790 ;
    END
  END w_mask_in[226]
  PIN w_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 108.790 0.460 109.250 ;
    END
  END w_mask_in[227]
  PIN w_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 109.250 0.460 109.710 ;
    END
  END w_mask_in[228]
  PIN w_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 109.710 0.460 110.170 ;
    END
  END w_mask_in[229]
  PIN w_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.170 0.460 110.630 ;
    END
  END w_mask_in[230]
  PIN w_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.630 0.460 111.090 ;
    END
  END w_mask_in[231]
  PIN w_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.090 0.460 111.550 ;
    END
  END w_mask_in[232]
  PIN w_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.550 0.460 112.010 ;
    END
  END w_mask_in[233]
  PIN w_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.010 0.460 112.470 ;
    END
  END w_mask_in[234]
  PIN w_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.470 0.460 112.930 ;
    END
  END w_mask_in[235]
  PIN w_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.930 0.460 113.390 ;
    END
  END w_mask_in[236]
  PIN w_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 113.390 0.460 113.850 ;
    END
  END w_mask_in[237]
  PIN w_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 113.850 0.460 114.310 ;
    END
  END w_mask_in[238]
  PIN w_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 114.310 0.460 114.770 ;
    END
  END w_mask_in[239]
  PIN w_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 114.770 0.460 115.230 ;
    END
  END w_mask_in[240]
  PIN w_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.230 0.460 115.690 ;
    END
  END w_mask_in[241]
  PIN w_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.690 0.460 116.150 ;
    END
  END w_mask_in[242]
  PIN w_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.150 0.460 116.610 ;
    END
  END w_mask_in[243]
  PIN w_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.610 0.460 117.070 ;
    END
  END w_mask_in[244]
  PIN w_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 117.070 0.460 117.530 ;
    END
  END w_mask_in[245]
  PIN w_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 117.530 0.460 117.990 ;
    END
  END w_mask_in[246]
  PIN w_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 117.990 0.460 118.450 ;
    END
  END w_mask_in[247]
  PIN w_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.450 0.460 118.910 ;
    END
  END w_mask_in[248]
  PIN w_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.910 0.460 119.370 ;
    END
  END w_mask_in[249]
  PIN w_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.370 0.460 119.830 ;
    END
  END w_mask_in[250]
  PIN w_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.830 0.460 120.290 ;
    END
  END w_mask_in[251]
  PIN w_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.290 0.460 120.750 ;
    END
  END w_mask_in[252]
  PIN w_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.750 0.460 121.210 ;
    END
  END w_mask_in[253]
  PIN w_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 121.210 0.460 121.670 ;
    END
  END w_mask_in[254]
  PIN w_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 121.670 0.460 122.130 ;
    END
  END w_mask_in[255]
  PIN w_mask_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 122.130 0.460 122.590 ;
    END
  END w_mask_in[256]
  PIN w_mask_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 122.590 0.460 123.050 ;
    END
  END w_mask_in[257]
  PIN w_mask_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.050 0.460 123.510 ;
    END
  END w_mask_in[258]
  PIN w_mask_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.510 0.460 123.970 ;
    END
  END w_mask_in[259]
  PIN w_mask_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.970 0.460 124.430 ;
    END
  END w_mask_in[260]
  PIN w_mask_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 124.430 0.460 124.890 ;
    END
  END w_mask_in[261]
  PIN w_mask_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 124.890 0.460 125.350 ;
    END
  END w_mask_in[262]
  PIN w_mask_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 125.350 0.460 125.810 ;
    END
  END w_mask_in[263]
  PIN w_mask_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 125.810 0.460 126.270 ;
    END
  END w_mask_in[264]
  PIN w_mask_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 126.270 0.460 126.730 ;
    END
  END w_mask_in[265]
  PIN w_mask_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 126.730 0.460 127.190 ;
    END
  END w_mask_in[266]
  PIN w_mask_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.190 0.460 127.650 ;
    END
  END w_mask_in[267]
  PIN w_mask_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.650 0.460 128.110 ;
    END
  END w_mask_in[268]
  PIN w_mask_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 128.110 0.460 128.570 ;
    END
  END w_mask_in[269]
  PIN w_mask_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 128.570 0.460 129.030 ;
    END
  END w_mask_in[270]
  PIN w_mask_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 129.030 0.460 129.490 ;
    END
  END w_mask_in[271]
  PIN w_mask_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 129.490 0.460 129.950 ;
    END
  END w_mask_in[272]
  PIN w_mask_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 129.950 0.460 130.410 ;
    END
  END w_mask_in[273]
  PIN w_mask_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.410 0.460 130.870 ;
    END
  END w_mask_in[274]
  PIN w_mask_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.870 0.460 131.330 ;
    END
  END w_mask_in[275]
  PIN w_mask_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.330 0.460 131.790 ;
    END
  END w_mask_in[276]
  PIN w_mask_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.790 0.460 132.250 ;
    END
  END w_mask_in[277]
  PIN w_mask_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 132.250 0.460 132.710 ;
    END
  END w_mask_in[278]
  PIN w_mask_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 132.710 0.460 133.170 ;
    END
  END w_mask_in[279]
  PIN w_mask_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.170 0.460 133.630 ;
    END
  END w_mask_in[280]
  PIN w_mask_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.630 0.460 134.090 ;
    END
  END w_mask_in[281]
  PIN w_mask_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.090 0.460 134.550 ;
    END
  END w_mask_in[282]
  PIN w_mask_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.550 0.460 135.010 ;
    END
  END w_mask_in[283]
  PIN w_mask_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.010 0.460 135.470 ;
    END
  END w_mask_in[284]
  PIN w_mask_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.470 0.460 135.930 ;
    END
  END w_mask_in[285]
  PIN w_mask_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.930 0.460 136.390 ;
    END
  END w_mask_in[286]
  PIN w_mask_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.390 0.460 136.850 ;
    END
  END w_mask_in[287]
  PIN w_mask_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.850 0.460 137.310 ;
    END
  END w_mask_in[288]
  PIN w_mask_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.310 0.460 137.770 ;
    END
  END w_mask_in[289]
  PIN w_mask_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.770 0.460 138.230 ;
    END
  END w_mask_in[290]
  PIN w_mask_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 138.230 0.460 138.690 ;
    END
  END w_mask_in[291]
  PIN w_mask_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 138.690 0.460 139.150 ;
    END
  END w_mask_in[292]
  PIN w_mask_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.150 0.460 139.610 ;
    END
  END w_mask_in[293]
  PIN w_mask_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.610 0.460 140.070 ;
    END
  END w_mask_in[294]
  PIN w_mask_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 140.070 0.460 140.530 ;
    END
  END w_mask_in[295]
  PIN w_mask_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 140.530 0.460 140.990 ;
    END
  END w_mask_in[296]
  PIN w_mask_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 140.990 0.460 141.450 ;
    END
  END w_mask_in[297]
  PIN w_mask_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.450 0.460 141.910 ;
    END
  END w_mask_in[298]
  PIN w_mask_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.910 0.460 142.370 ;
    END
  END w_mask_in[299]
  PIN w_mask_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.370 0.460 142.830 ;
    END
  END w_mask_in[300]
  PIN w_mask_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.830 0.460 143.290 ;
    END
  END w_mask_in[301]
  PIN w_mask_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.290 0.460 143.750 ;
    END
  END w_mask_in[302]
  PIN w_mask_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.750 0.460 144.210 ;
    END
  END w_mask_in[303]
  PIN w_mask_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.210 0.460 144.670 ;
    END
  END w_mask_in[304]
  PIN w_mask_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.670 0.460 145.130 ;
    END
  END w_mask_in[305]
  PIN w_mask_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.130 0.460 145.590 ;
    END
  END w_mask_in[306]
  PIN w_mask_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.590 0.460 146.050 ;
    END
  END w_mask_in[307]
  PIN w_mask_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.050 0.460 146.510 ;
    END
  END w_mask_in[308]
  PIN w_mask_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.510 0.460 146.970 ;
    END
  END w_mask_in[309]
  PIN w_mask_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.970 0.460 147.430 ;
    END
  END w_mask_in[310]
  PIN w_mask_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 147.430 0.460 147.890 ;
    END
  END w_mask_in[311]
  PIN w_mask_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 147.890 0.460 148.350 ;
    END
  END w_mask_in[312]
  PIN w_mask_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.350 0.460 148.810 ;
    END
  END w_mask_in[313]
  PIN w_mask_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.810 0.460 149.270 ;
    END
  END w_mask_in[314]
  PIN w_mask_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.270 0.460 149.730 ;
    END
  END w_mask_in[315]
  PIN w_mask_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.730 0.460 150.190 ;
    END
  END w_mask_in[316]
  PIN w_mask_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.190 0.460 150.650 ;
    END
  END w_mask_in[317]
  PIN w_mask_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.650 0.460 151.110 ;
    END
  END w_mask_in[318]
  PIN w_mask_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.110 0.460 151.570 ;
    END
  END w_mask_in[319]
  PIN w_mask_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.570 0.460 152.030 ;
    END
  END w_mask_in[320]
  PIN w_mask_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.030 0.460 152.490 ;
    END
  END w_mask_in[321]
  PIN w_mask_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.490 0.460 152.950 ;
    END
  END w_mask_in[322]
  PIN w_mask_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.950 0.460 153.410 ;
    END
  END w_mask_in[323]
  PIN w_mask_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.410 0.460 153.870 ;
    END
  END w_mask_in[324]
  PIN w_mask_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.870 0.460 154.330 ;
    END
  END w_mask_in[325]
  PIN w_mask_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.330 0.460 154.790 ;
    END
  END w_mask_in[326]
  PIN w_mask_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.790 0.460 155.250 ;
    END
  END w_mask_in[327]
  PIN w_mask_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 155.250 0.460 155.710 ;
    END
  END w_mask_in[328]
  PIN w_mask_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 155.710 0.460 156.170 ;
    END
  END w_mask_in[329]
  PIN w_mask_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.170 0.460 156.630 ;
    END
  END w_mask_in[330]
  PIN w_mask_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.630 0.460 157.090 ;
    END
  END w_mask_in[331]
  PIN w_mask_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.090 0.460 157.550 ;
    END
  END w_mask_in[332]
  PIN w_mask_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.550 0.460 158.010 ;
    END
  END w_mask_in[333]
  PIN w_mask_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.010 0.460 158.470 ;
    END
  END w_mask_in[334]
  PIN w_mask_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.470 0.460 158.930 ;
    END
  END w_mask_in[335]
  PIN w_mask_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.930 0.460 159.390 ;
    END
  END w_mask_in[336]
  PIN w_mask_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 159.390 0.460 159.850 ;
    END
  END w_mask_in[337]
  PIN w_mask_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 159.850 0.460 160.310 ;
    END
  END w_mask_in[338]
  PIN w_mask_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 160.310 0.460 160.770 ;
    END
  END w_mask_in[339]
  PIN w_mask_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 160.770 0.460 161.230 ;
    END
  END w_mask_in[340]
  PIN w_mask_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.230 0.460 161.690 ;
    END
  END w_mask_in[341]
  PIN w_mask_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.690 0.460 162.150 ;
    END
  END w_mask_in[342]
  PIN w_mask_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.150 0.460 162.610 ;
    END
  END w_mask_in[343]
  PIN w_mask_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.610 0.460 163.070 ;
    END
  END w_mask_in[344]
  PIN w_mask_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.070 0.460 163.530 ;
    END
  END w_mask_in[345]
  PIN w_mask_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.530 0.460 163.990 ;
    END
  END w_mask_in[346]
  PIN w_mask_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.990 0.460 164.450 ;
    END
  END w_mask_in[347]
  PIN w_mask_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.450 0.460 164.910 ;
    END
  END w_mask_in[348]
  PIN w_mask_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.910 0.460 165.370 ;
    END
  END w_mask_in[349]
  PIN w_mask_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.370 0.460 165.830 ;
    END
  END w_mask_in[350]
  PIN w_mask_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.830 0.460 166.290 ;
    END
  END w_mask_in[351]
  PIN w_mask_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.290 0.460 166.750 ;
    END
  END w_mask_in[352]
  PIN w_mask_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.750 0.460 167.210 ;
    END
  END w_mask_in[353]
  PIN w_mask_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.210 0.460 167.670 ;
    END
  END w_mask_in[354]
  PIN w_mask_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.670 0.460 168.130 ;
    END
  END w_mask_in[355]
  PIN w_mask_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.130 0.460 168.590 ;
    END
  END w_mask_in[356]
  PIN w_mask_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.590 0.460 169.050 ;
    END
  END w_mask_in[357]
  PIN w_mask_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.050 0.460 169.510 ;
    END
  END w_mask_in[358]
  PIN w_mask_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.510 0.460 169.970 ;
    END
  END w_mask_in[359]
  PIN w_mask_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.970 0.460 170.430 ;
    END
  END w_mask_in[360]
  PIN w_mask_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 170.430 0.460 170.890 ;
    END
  END w_mask_in[361]
  PIN w_mask_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 170.890 0.460 171.350 ;
    END
  END w_mask_in[362]
  PIN w_mask_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 171.350 0.460 171.810 ;
    END
  END w_mask_in[363]
  PIN w_mask_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 171.810 0.460 172.270 ;
    END
  END w_mask_in[364]
  PIN w_mask_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 172.270 0.460 172.730 ;
    END
  END w_mask_in[365]
  PIN w_mask_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 172.730 0.460 173.190 ;
    END
  END w_mask_in[366]
  PIN w_mask_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 173.190 0.460 173.650 ;
    END
  END w_mask_in[367]
  PIN w_mask_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 173.650 0.460 174.110 ;
    END
  END w_mask_in[368]
  PIN w_mask_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 174.110 0.460 174.570 ;
    END
  END w_mask_in[369]
  PIN w_mask_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 174.570 0.460 175.030 ;
    END
  END w_mask_in[370]
  PIN w_mask_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.030 0.460 175.490 ;
    END
  END w_mask_in[371]
  PIN w_mask_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.490 0.460 175.950 ;
    END
  END w_mask_in[372]
  PIN w_mask_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.950 0.460 176.410 ;
    END
  END w_mask_in[373]
  PIN w_mask_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 176.410 0.460 176.870 ;
    END
  END w_mask_in[374]
  PIN w_mask_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 176.870 0.460 177.330 ;
    END
  END w_mask_in[375]
  PIN w_mask_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 177.330 0.460 177.790 ;
    END
  END w_mask_in[376]
  PIN w_mask_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 177.790 0.460 178.250 ;
    END
  END w_mask_in[377]
  PIN w_mask_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 178.250 0.460 178.710 ;
    END
  END w_mask_in[378]
  PIN w_mask_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 178.710 0.460 179.170 ;
    END
  END w_mask_in[379]
  PIN w_mask_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 179.170 0.460 179.630 ;
    END
  END w_mask_in[380]
  PIN w_mask_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 179.630 0.460 180.090 ;
    END
  END w_mask_in[381]
  PIN w_mask_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 180.090 0.460 180.550 ;
    END
  END w_mask_in[382]
  PIN w_mask_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 180.550 0.460 181.010 ;
    END
  END w_mask_in[383]
  PIN w_mask_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 181.010 0.460 181.470 ;
    END
  END w_mask_in[384]
  PIN w_mask_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 181.470 0.460 181.930 ;
    END
  END w_mask_in[385]
  PIN w_mask_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 181.930 0.460 182.390 ;
    END
  END w_mask_in[386]
  PIN w_mask_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 182.390 0.460 182.850 ;
    END
  END w_mask_in[387]
  PIN w_mask_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 182.850 0.460 183.310 ;
    END
  END w_mask_in[388]
  PIN w_mask_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 183.310 0.460 183.770 ;
    END
  END w_mask_in[389]
  PIN w_mask_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 183.770 0.460 184.230 ;
    END
  END w_mask_in[390]
  PIN w_mask_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 184.230 0.460 184.690 ;
    END
  END w_mask_in[391]
  PIN w_mask_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 184.690 0.460 185.150 ;
    END
  END w_mask_in[392]
  PIN w_mask_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 185.150 0.460 185.610 ;
    END
  END w_mask_in[393]
  PIN w_mask_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 185.610 0.460 186.070 ;
    END
  END w_mask_in[394]
  PIN w_mask_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.070 0.460 186.530 ;
    END
  END w_mask_in[395]
  PIN w_mask_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.530 0.460 186.990 ;
    END
  END w_mask_in[396]
  PIN w_mask_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.990 0.460 187.450 ;
    END
  END w_mask_in[397]
  PIN w_mask_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 187.450 0.460 187.910 ;
    END
  END w_mask_in[398]
  PIN w_mask_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 187.910 0.460 188.370 ;
    END
  END w_mask_in[399]
  PIN w_mask_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 188.370 0.460 188.830 ;
    END
  END w_mask_in[400]
  PIN w_mask_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 188.830 0.460 189.290 ;
    END
  END w_mask_in[401]
  PIN w_mask_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 189.290 0.460 189.750 ;
    END
  END w_mask_in[402]
  PIN w_mask_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 189.750 0.460 190.210 ;
    END
  END w_mask_in[403]
  PIN w_mask_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 190.210 0.460 190.670 ;
    END
  END w_mask_in[404]
  PIN w_mask_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 190.670 0.460 191.130 ;
    END
  END w_mask_in[405]
  PIN w_mask_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 191.130 0.460 191.590 ;
    END
  END w_mask_in[406]
  PIN w_mask_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 191.590 0.460 192.050 ;
    END
  END w_mask_in[407]
  PIN w_mask_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 192.050 0.460 192.510 ;
    END
  END w_mask_in[408]
  PIN w_mask_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 192.510 0.460 192.970 ;
    END
  END w_mask_in[409]
  PIN w_mask_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 192.970 0.460 193.430 ;
    END
  END w_mask_in[410]
  PIN w_mask_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 193.430 0.460 193.890 ;
    END
  END w_mask_in[411]
  PIN w_mask_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 193.890 0.460 194.350 ;
    END
  END w_mask_in[412]
  PIN w_mask_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.350 0.460 194.810 ;
    END
  END w_mask_in[413]
  PIN w_mask_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.810 0.460 195.270 ;
    END
  END w_mask_in[414]
  PIN w_mask_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.270 0.460 195.730 ;
    END
  END w_mask_in[415]
  PIN w_mask_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.730 0.460 196.190 ;
    END
  END w_mask_in[416]
  PIN w_mask_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 196.190 0.460 196.650 ;
    END
  END w_mask_in[417]
  PIN w_mask_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 196.650 0.460 197.110 ;
    END
  END w_mask_in[418]
  PIN w_mask_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 197.110 0.460 197.570 ;
    END
  END w_mask_in[419]
  PIN w_mask_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 197.570 0.460 198.030 ;
    END
  END w_mask_in[420]
  PIN w_mask_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 198.030 0.460 198.490 ;
    END
  END w_mask_in[421]
  PIN w_mask_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 198.490 0.460 198.950 ;
    END
  END w_mask_in[422]
  PIN w_mask_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 198.950 0.460 199.410 ;
    END
  END w_mask_in[423]
  PIN w_mask_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 199.410 0.460 199.870 ;
    END
  END w_mask_in[424]
  PIN w_mask_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 199.870 0.460 200.330 ;
    END
  END w_mask_in[425]
  PIN w_mask_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 200.330 0.460 200.790 ;
    END
  END w_mask_in[426]
  PIN w_mask_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 200.790 0.460 201.250 ;
    END
  END w_mask_in[427]
  PIN w_mask_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 201.250 0.460 201.710 ;
    END
  END w_mask_in[428]
  PIN w_mask_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 201.710 0.460 202.170 ;
    END
  END w_mask_in[429]
  PIN w_mask_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 202.170 0.460 202.630 ;
    END
  END w_mask_in[430]
  PIN w_mask_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 202.630 0.460 203.090 ;
    END
  END w_mask_in[431]
  PIN w_mask_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 203.090 0.460 203.550 ;
    END
  END w_mask_in[432]
  PIN w_mask_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 203.550 0.460 204.010 ;
    END
  END w_mask_in[433]
  PIN w_mask_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 204.010 0.460 204.470 ;
    END
  END w_mask_in[434]
  PIN w_mask_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 204.470 0.460 204.930 ;
    END
  END w_mask_in[435]
  PIN w_mask_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 204.930 0.460 205.390 ;
    END
  END w_mask_in[436]
  PIN w_mask_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.390 0.460 205.850 ;
    END
  END w_mask_in[437]
  PIN w_mask_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.850 0.460 206.310 ;
    END
  END w_mask_in[438]
  PIN w_mask_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 206.310 0.460 206.770 ;
    END
  END w_mask_in[439]
  PIN w_mask_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 206.770 0.460 207.230 ;
    END
  END w_mask_in[440]
  PIN w_mask_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 207.230 0.460 207.690 ;
    END
  END w_mask_in[441]
  PIN w_mask_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 207.690 0.460 208.150 ;
    END
  END w_mask_in[442]
  PIN w_mask_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 208.150 0.460 208.610 ;
    END
  END w_mask_in[443]
  PIN w_mask_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 208.610 0.460 209.070 ;
    END
  END w_mask_in[444]
  PIN w_mask_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.070 0.460 209.530 ;
    END
  END w_mask_in[445]
  PIN w_mask_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.530 0.460 209.990 ;
    END
  END w_mask_in[446]
  PIN w_mask_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.990 0.460 210.450 ;
    END
  END w_mask_in[447]
  PIN w_mask_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 210.450 0.460 210.910 ;
    END
  END w_mask_in[448]
  PIN w_mask_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 210.910 0.460 211.370 ;
    END
  END w_mask_in[449]
  PIN w_mask_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 211.370 0.460 211.830 ;
    END
  END w_mask_in[450]
  PIN w_mask_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 211.830 0.460 212.290 ;
    END
  END w_mask_in[451]
  PIN w_mask_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 212.290 0.460 212.750 ;
    END
  END w_mask_in[452]
  PIN w_mask_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 212.750 0.460 213.210 ;
    END
  END w_mask_in[453]
  PIN w_mask_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 213.210 0.460 213.670 ;
    END
  END w_mask_in[454]
  PIN w_mask_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 213.670 0.460 214.130 ;
    END
  END w_mask_in[455]
  PIN w_mask_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 214.130 0.460 214.590 ;
    END
  END w_mask_in[456]
  PIN w_mask_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 214.590 0.460 215.050 ;
    END
  END w_mask_in[457]
  PIN w_mask_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 215.050 0.460 215.510 ;
    END
  END w_mask_in[458]
  PIN w_mask_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 215.510 0.460 215.970 ;
    END
  END w_mask_in[459]
  PIN w_mask_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 215.970 0.460 216.430 ;
    END
  END w_mask_in[460]
  PIN w_mask_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.430 0.460 216.890 ;
    END
  END w_mask_in[461]
  PIN w_mask_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.890 0.460 217.350 ;
    END
  END w_mask_in[462]
  PIN w_mask_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 217.350 0.460 217.810 ;
    END
  END w_mask_in[463]
  PIN w_mask_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 217.810 0.460 218.270 ;
    END
  END w_mask_in[464]
  PIN w_mask_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 218.270 0.460 218.730 ;
    END
  END w_mask_in[465]
  PIN w_mask_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 218.730 0.460 219.190 ;
    END
  END w_mask_in[466]
  PIN w_mask_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 219.190 0.460 219.650 ;
    END
  END w_mask_in[467]
  PIN w_mask_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 219.650 0.460 220.110 ;
    END
  END w_mask_in[468]
  PIN w_mask_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.110 0.460 220.570 ;
    END
  END w_mask_in[469]
  PIN w_mask_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.570 0.460 221.030 ;
    END
  END w_mask_in[470]
  PIN w_mask_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 221.030 0.460 221.490 ;
    END
  END w_mask_in[471]
  PIN w_mask_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 221.490 0.460 221.950 ;
    END
  END w_mask_in[472]
  PIN w_mask_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 221.950 0.460 222.410 ;
    END
  END w_mask_in[473]
  PIN w_mask_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 222.410 0.460 222.870 ;
    END
  END w_mask_in[474]
  PIN w_mask_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 222.870 0.460 223.330 ;
    END
  END w_mask_in[475]
  PIN w_mask_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.330 0.460 223.790 ;
    END
  END w_mask_in[476]
  PIN w_mask_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.790 0.460 224.250 ;
    END
  END w_mask_in[477]
  PIN w_mask_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 224.250 0.460 224.710 ;
    END
  END w_mask_in[478]
  PIN w_mask_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 224.710 0.460 225.170 ;
    END
  END w_mask_in[479]
  PIN w_mask_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 225.170 0.460 225.630 ;
    END
  END w_mask_in[480]
  PIN w_mask_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 225.630 0.460 226.090 ;
    END
  END w_mask_in[481]
  PIN w_mask_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 226.090 0.460 226.550 ;
    END
  END w_mask_in[482]
  PIN w_mask_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 226.550 0.460 227.010 ;
    END
  END w_mask_in[483]
  PIN w_mask_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 227.010 0.460 227.470 ;
    END
  END w_mask_in[484]
  PIN w_mask_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 227.470 0.460 227.930 ;
    END
  END w_mask_in[485]
  PIN w_mask_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 227.930 0.460 228.390 ;
    END
  END w_mask_in[486]
  PIN w_mask_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 228.390 0.460 228.850 ;
    END
  END w_mask_in[487]
  PIN w_mask_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 228.850 0.460 229.310 ;
    END
  END w_mask_in[488]
  PIN w_mask_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 229.310 0.460 229.770 ;
    END
  END w_mask_in[489]
  PIN w_mask_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 229.770 0.460 230.230 ;
    END
  END w_mask_in[490]
  PIN w_mask_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 230.230 0.460 230.690 ;
    END
  END w_mask_in[491]
  PIN w_mask_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 230.690 0.460 231.150 ;
    END
  END w_mask_in[492]
  PIN w_mask_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 231.150 0.460 231.610 ;
    END
  END w_mask_in[493]
  PIN w_mask_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 231.610 0.460 232.070 ;
    END
  END w_mask_in[494]
  PIN w_mask_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 232.070 0.460 232.530 ;
    END
  END w_mask_in[495]
  PIN w_mask_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 232.530 0.460 232.990 ;
    END
  END w_mask_in[496]
  PIN w_mask_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 232.990 0.460 233.450 ;
    END
  END w_mask_in[497]
  PIN w_mask_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 233.450 0.460 233.910 ;
    END
  END w_mask_in[498]
  PIN w_mask_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 233.910 0.460 234.370 ;
    END
  END w_mask_in[499]
  PIN w_mask_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 234.370 0.460 234.830 ;
    END
  END w_mask_in[500]
  PIN w_mask_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 234.830 0.460 235.290 ;
    END
  END w_mask_in[501]
  PIN w_mask_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 235.290 0.460 235.750 ;
    END
  END w_mask_in[502]
  PIN w_mask_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 235.750 0.460 236.210 ;
    END
  END w_mask_in[503]
  PIN w_mask_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 236.210 0.460 236.670 ;
    END
  END w_mask_in[504]
  PIN w_mask_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 236.670 0.460 237.130 ;
    END
  END w_mask_in[505]
  PIN w_mask_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 237.130 0.460 237.590 ;
    END
  END w_mask_in[506]
  PIN w_mask_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 237.590 0.460 238.050 ;
    END
  END w_mask_in[507]
  PIN w_mask_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 238.050 0.460 238.510 ;
    END
  END w_mask_in[508]
  PIN w_mask_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 238.510 0.460 238.970 ;
    END
  END w_mask_in[509]
  PIN w_mask_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 238.970 0.460 239.430 ;
    END
  END w_mask_in[510]
  PIN w_mask_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 239.430 0.460 239.890 ;
    END
  END w_mask_in[511]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 322.230 0.460 322.690 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 322.690 0.460 323.150 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 323.150 0.460 323.610 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 323.610 0.460 324.070 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 324.070 0.460 324.530 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 324.530 0.460 324.990 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 324.990 0.460 325.450 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 325.450 0.460 325.910 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 325.910 0.460 326.370 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 326.370 0.460 326.830 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 326.830 0.460 327.290 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.290 0.460 327.750 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.750 0.460 328.210 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 328.210 0.460 328.670 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 328.670 0.460 329.130 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 329.130 0.460 329.590 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 329.590 0.460 330.050 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.050 0.460 330.510 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.510 0.460 330.970 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.970 0.460 331.430 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 331.430 0.460 331.890 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 331.890 0.460 332.350 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 332.350 0.460 332.810 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 332.810 0.460 333.270 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.270 0.460 333.730 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.730 0.460 334.190 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 334.190 0.460 334.650 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 334.650 0.460 335.110 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 335.110 0.460 335.570 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 335.570 0.460 336.030 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 336.030 0.460 336.490 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 336.490 0.460 336.950 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 336.950 0.460 337.410 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.410 0.460 337.870 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.870 0.460 338.330 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 338.330 0.460 338.790 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 338.790 0.460 339.250 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 339.250 0.460 339.710 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 339.710 0.460 340.170 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 340.170 0.460 340.630 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 340.630 0.460 341.090 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 341.090 0.460 341.550 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 341.550 0.460 342.010 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 342.010 0.460 342.470 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 342.470 0.460 342.930 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 342.930 0.460 343.390 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 343.390 0.460 343.850 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 343.850 0.460 344.310 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 344.310 0.460 344.770 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 344.770 0.460 345.230 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 345.230 0.460 345.690 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 345.690 0.460 346.150 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 346.150 0.460 346.610 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 346.610 0.460 347.070 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 347.070 0.460 347.530 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 347.530 0.460 347.990 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 347.990 0.460 348.450 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 348.450 0.460 348.910 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 348.910 0.460 349.370 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 349.370 0.460 349.830 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 349.830 0.460 350.290 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 350.290 0.460 350.750 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 350.750 0.460 351.210 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 351.210 0.460 351.670 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 351.670 0.460 352.130 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 352.130 0.460 352.590 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 352.590 0.460 353.050 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 353.050 0.460 353.510 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 353.510 0.460 353.970 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 353.970 0.460 354.430 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 354.430 0.460 354.890 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 354.890 0.460 355.350 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 355.350 0.460 355.810 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 355.810 0.460 356.270 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 356.270 0.460 356.730 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 356.730 0.460 357.190 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 357.190 0.460 357.650 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 357.650 0.460 358.110 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 358.110 0.460 358.570 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 358.570 0.460 359.030 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 359.030 0.460 359.490 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 359.490 0.460 359.950 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 359.950 0.460 360.410 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 360.410 0.460 360.870 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 360.870 0.460 361.330 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 361.330 0.460 361.790 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 361.790 0.460 362.250 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 362.250 0.460 362.710 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 362.710 0.460 363.170 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 363.170 0.460 363.630 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 363.630 0.460 364.090 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 364.090 0.460 364.550 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 364.550 0.460 365.010 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 365.010 0.460 365.470 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 365.470 0.460 365.930 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 365.930 0.460 366.390 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 366.390 0.460 366.850 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 366.850 0.460 367.310 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 367.310 0.460 367.770 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 367.770 0.460 368.230 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 368.230 0.460 368.690 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 368.690 0.460 369.150 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 369.150 0.460 369.610 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 369.610 0.460 370.070 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 370.070 0.460 370.530 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 370.530 0.460 370.990 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 370.990 0.460 371.450 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 371.450 0.460 371.910 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 371.910 0.460 372.370 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 372.370 0.460 372.830 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 372.830 0.460 373.290 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 373.290 0.460 373.750 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 373.750 0.460 374.210 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 374.210 0.460 374.670 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 374.670 0.460 375.130 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 375.130 0.460 375.590 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 375.590 0.460 376.050 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 376.050 0.460 376.510 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 376.510 0.460 376.970 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 376.970 0.460 377.430 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 377.430 0.460 377.890 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 377.890 0.460 378.350 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 378.350 0.460 378.810 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 378.810 0.460 379.270 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 379.270 0.460 379.730 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 379.730 0.460 380.190 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 380.190 0.460 380.650 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 380.650 0.460 381.110 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 381.110 0.460 381.570 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 381.570 0.460 382.030 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 382.030 0.460 382.490 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 382.490 0.460 382.950 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 382.950 0.460 383.410 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 383.410 0.460 383.870 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 383.870 0.460 384.330 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 384.330 0.460 384.790 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 384.790 0.460 385.250 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 385.250 0.460 385.710 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 385.710 0.460 386.170 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 386.170 0.460 386.630 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 386.630 0.460 387.090 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 387.090 0.460 387.550 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 387.550 0.460 388.010 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 388.010 0.460 388.470 ;
    END
  END rd_out[143]
  PIN rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 388.470 0.460 388.930 ;
    END
  END rd_out[144]
  PIN rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 388.930 0.460 389.390 ;
    END
  END rd_out[145]
  PIN rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 389.390 0.460 389.850 ;
    END
  END rd_out[146]
  PIN rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 389.850 0.460 390.310 ;
    END
  END rd_out[147]
  PIN rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 390.310 0.460 390.770 ;
    END
  END rd_out[148]
  PIN rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 390.770 0.460 391.230 ;
    END
  END rd_out[149]
  PIN rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 391.230 0.460 391.690 ;
    END
  END rd_out[150]
  PIN rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 391.690 0.460 392.150 ;
    END
  END rd_out[151]
  PIN rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 392.150 0.460 392.610 ;
    END
  END rd_out[152]
  PIN rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 392.610 0.460 393.070 ;
    END
  END rd_out[153]
  PIN rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 393.070 0.460 393.530 ;
    END
  END rd_out[154]
  PIN rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 393.530 0.460 393.990 ;
    END
  END rd_out[155]
  PIN rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 393.990 0.460 394.450 ;
    END
  END rd_out[156]
  PIN rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 394.450 0.460 394.910 ;
    END
  END rd_out[157]
  PIN rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 394.910 0.460 395.370 ;
    END
  END rd_out[158]
  PIN rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 395.370 0.460 395.830 ;
    END
  END rd_out[159]
  PIN rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 395.830 0.460 396.290 ;
    END
  END rd_out[160]
  PIN rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 396.290 0.460 396.750 ;
    END
  END rd_out[161]
  PIN rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 396.750 0.460 397.210 ;
    END
  END rd_out[162]
  PIN rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 397.210 0.460 397.670 ;
    END
  END rd_out[163]
  PIN rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 397.670 0.460 398.130 ;
    END
  END rd_out[164]
  PIN rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 398.130 0.460 398.590 ;
    END
  END rd_out[165]
  PIN rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 398.590 0.460 399.050 ;
    END
  END rd_out[166]
  PIN rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.050 0.460 399.510 ;
    END
  END rd_out[167]
  PIN rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.510 0.460 399.970 ;
    END
  END rd_out[168]
  PIN rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.970 0.460 400.430 ;
    END
  END rd_out[169]
  PIN rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 400.430 0.460 400.890 ;
    END
  END rd_out[170]
  PIN rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 400.890 0.460 401.350 ;
    END
  END rd_out[171]
  PIN rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 401.350 0.460 401.810 ;
    END
  END rd_out[172]
  PIN rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 401.810 0.460 402.270 ;
    END
  END rd_out[173]
  PIN rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 402.270 0.460 402.730 ;
    END
  END rd_out[174]
  PIN rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 402.730 0.460 403.190 ;
    END
  END rd_out[175]
  PIN rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 403.190 0.460 403.650 ;
    END
  END rd_out[176]
  PIN rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 403.650 0.460 404.110 ;
    END
  END rd_out[177]
  PIN rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 404.110 0.460 404.570 ;
    END
  END rd_out[178]
  PIN rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 404.570 0.460 405.030 ;
    END
  END rd_out[179]
  PIN rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 405.030 0.460 405.490 ;
    END
  END rd_out[180]
  PIN rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 405.490 0.460 405.950 ;
    END
  END rd_out[181]
  PIN rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 405.950 0.460 406.410 ;
    END
  END rd_out[182]
  PIN rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 406.410 0.460 406.870 ;
    END
  END rd_out[183]
  PIN rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 406.870 0.460 407.330 ;
    END
  END rd_out[184]
  PIN rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 407.330 0.460 407.790 ;
    END
  END rd_out[185]
  PIN rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 407.790 0.460 408.250 ;
    END
  END rd_out[186]
  PIN rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 408.250 0.460 408.710 ;
    END
  END rd_out[187]
  PIN rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 408.710 0.460 409.170 ;
    END
  END rd_out[188]
  PIN rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.170 0.460 409.630 ;
    END
  END rd_out[189]
  PIN rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.630 0.460 410.090 ;
    END
  END rd_out[190]
  PIN rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 410.090 0.460 410.550 ;
    END
  END rd_out[191]
  PIN rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 410.550 0.460 411.010 ;
    END
  END rd_out[192]
  PIN rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 411.010 0.460 411.470 ;
    END
  END rd_out[193]
  PIN rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 411.470 0.460 411.930 ;
    END
  END rd_out[194]
  PIN rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 411.930 0.460 412.390 ;
    END
  END rd_out[195]
  PIN rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 412.390 0.460 412.850 ;
    END
  END rd_out[196]
  PIN rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 412.850 0.460 413.310 ;
    END
  END rd_out[197]
  PIN rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 413.310 0.460 413.770 ;
    END
  END rd_out[198]
  PIN rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 413.770 0.460 414.230 ;
    END
  END rd_out[199]
  PIN rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 414.230 0.460 414.690 ;
    END
  END rd_out[200]
  PIN rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 414.690 0.460 415.150 ;
    END
  END rd_out[201]
  PIN rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 415.150 0.460 415.610 ;
    END
  END rd_out[202]
  PIN rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 415.610 0.460 416.070 ;
    END
  END rd_out[203]
  PIN rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 416.070 0.460 416.530 ;
    END
  END rd_out[204]
  PIN rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 416.530 0.460 416.990 ;
    END
  END rd_out[205]
  PIN rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 416.990 0.460 417.450 ;
    END
  END rd_out[206]
  PIN rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 417.450 0.460 417.910 ;
    END
  END rd_out[207]
  PIN rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 417.910 0.460 418.370 ;
    END
  END rd_out[208]
  PIN rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 418.370 0.460 418.830 ;
    END
  END rd_out[209]
  PIN rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 418.830 0.460 419.290 ;
    END
  END rd_out[210]
  PIN rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 419.290 0.460 419.750 ;
    END
  END rd_out[211]
  PIN rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 419.750 0.460 420.210 ;
    END
  END rd_out[212]
  PIN rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 420.210 0.460 420.670 ;
    END
  END rd_out[213]
  PIN rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 420.670 0.460 421.130 ;
    END
  END rd_out[214]
  PIN rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 421.130 0.460 421.590 ;
    END
  END rd_out[215]
  PIN rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 421.590 0.460 422.050 ;
    END
  END rd_out[216]
  PIN rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 422.050 0.460 422.510 ;
    END
  END rd_out[217]
  PIN rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 422.510 0.460 422.970 ;
    END
  END rd_out[218]
  PIN rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 422.970 0.460 423.430 ;
    END
  END rd_out[219]
  PIN rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 423.430 0.460 423.890 ;
    END
  END rd_out[220]
  PIN rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 423.890 0.460 424.350 ;
    END
  END rd_out[221]
  PIN rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 424.350 0.460 424.810 ;
    END
  END rd_out[222]
  PIN rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 424.810 0.460 425.270 ;
    END
  END rd_out[223]
  PIN rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 425.270 0.460 425.730 ;
    END
  END rd_out[224]
  PIN rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 425.730 0.460 426.190 ;
    END
  END rd_out[225]
  PIN rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 426.190 0.460 426.650 ;
    END
  END rd_out[226]
  PIN rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 426.650 0.460 427.110 ;
    END
  END rd_out[227]
  PIN rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 427.110 0.460 427.570 ;
    END
  END rd_out[228]
  PIN rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 427.570 0.460 428.030 ;
    END
  END rd_out[229]
  PIN rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 428.030 0.460 428.490 ;
    END
  END rd_out[230]
  PIN rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 428.490 0.460 428.950 ;
    END
  END rd_out[231]
  PIN rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 428.950 0.460 429.410 ;
    END
  END rd_out[232]
  PIN rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 429.410 0.460 429.870 ;
    END
  END rd_out[233]
  PIN rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 429.870 0.460 430.330 ;
    END
  END rd_out[234]
  PIN rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 430.330 0.460 430.790 ;
    END
  END rd_out[235]
  PIN rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 430.790 0.460 431.250 ;
    END
  END rd_out[236]
  PIN rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 431.250 0.460 431.710 ;
    END
  END rd_out[237]
  PIN rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 431.710 0.460 432.170 ;
    END
  END rd_out[238]
  PIN rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 432.170 0.460 432.630 ;
    END
  END rd_out[239]
  PIN rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 432.630 0.460 433.090 ;
    END
  END rd_out[240]
  PIN rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 433.090 0.460 433.550 ;
    END
  END rd_out[241]
  PIN rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 433.550 0.460 434.010 ;
    END
  END rd_out[242]
  PIN rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 434.010 0.460 434.470 ;
    END
  END rd_out[243]
  PIN rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 434.470 0.460 434.930 ;
    END
  END rd_out[244]
  PIN rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 434.930 0.460 435.390 ;
    END
  END rd_out[245]
  PIN rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 435.390 0.460 435.850 ;
    END
  END rd_out[246]
  PIN rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 435.850 0.460 436.310 ;
    END
  END rd_out[247]
  PIN rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 436.310 0.460 436.770 ;
    END
  END rd_out[248]
  PIN rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 436.770 0.460 437.230 ;
    END
  END rd_out[249]
  PIN rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 437.230 0.460 437.690 ;
    END
  END rd_out[250]
  PIN rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 437.690 0.460 438.150 ;
    END
  END rd_out[251]
  PIN rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 438.150 0.460 438.610 ;
    END
  END rd_out[252]
  PIN rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 438.610 0.460 439.070 ;
    END
  END rd_out[253]
  PIN rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 439.070 0.460 439.530 ;
    END
  END rd_out[254]
  PIN rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 439.530 0.460 439.990 ;
    END
  END rd_out[255]
  PIN rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 439.990 0.460 440.450 ;
    END
  END rd_out[256]
  PIN rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 440.450 0.460 440.910 ;
    END
  END rd_out[257]
  PIN rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 440.910 0.460 441.370 ;
    END
  END rd_out[258]
  PIN rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 441.370 0.460 441.830 ;
    END
  END rd_out[259]
  PIN rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 441.830 0.460 442.290 ;
    END
  END rd_out[260]
  PIN rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 442.290 0.460 442.750 ;
    END
  END rd_out[261]
  PIN rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 442.750 0.460 443.210 ;
    END
  END rd_out[262]
  PIN rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 443.210 0.460 443.670 ;
    END
  END rd_out[263]
  PIN rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 443.670 0.460 444.130 ;
    END
  END rd_out[264]
  PIN rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 444.130 0.460 444.590 ;
    END
  END rd_out[265]
  PIN rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 444.590 0.460 445.050 ;
    END
  END rd_out[266]
  PIN rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 445.050 0.460 445.510 ;
    END
  END rd_out[267]
  PIN rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 445.510 0.460 445.970 ;
    END
  END rd_out[268]
  PIN rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 445.970 0.460 446.430 ;
    END
  END rd_out[269]
  PIN rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 446.430 0.460 446.890 ;
    END
  END rd_out[270]
  PIN rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 446.890 0.460 447.350 ;
    END
  END rd_out[271]
  PIN rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 447.350 0.460 447.810 ;
    END
  END rd_out[272]
  PIN rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 447.810 0.460 448.270 ;
    END
  END rd_out[273]
  PIN rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 448.270 0.460 448.730 ;
    END
  END rd_out[274]
  PIN rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 448.730 0.460 449.190 ;
    END
  END rd_out[275]
  PIN rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 449.190 0.460 449.650 ;
    END
  END rd_out[276]
  PIN rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 449.650 0.460 450.110 ;
    END
  END rd_out[277]
  PIN rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 450.110 0.460 450.570 ;
    END
  END rd_out[278]
  PIN rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 450.570 0.460 451.030 ;
    END
  END rd_out[279]
  PIN rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 451.030 0.460 451.490 ;
    END
  END rd_out[280]
  PIN rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 451.490 0.460 451.950 ;
    END
  END rd_out[281]
  PIN rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 451.950 0.460 452.410 ;
    END
  END rd_out[282]
  PIN rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 452.410 0.460 452.870 ;
    END
  END rd_out[283]
  PIN rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 452.870 0.460 453.330 ;
    END
  END rd_out[284]
  PIN rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 453.330 0.460 453.790 ;
    END
  END rd_out[285]
  PIN rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 453.790 0.460 454.250 ;
    END
  END rd_out[286]
  PIN rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 454.250 0.460 454.710 ;
    END
  END rd_out[287]
  PIN rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 454.710 0.460 455.170 ;
    END
  END rd_out[288]
  PIN rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 455.170 0.460 455.630 ;
    END
  END rd_out[289]
  PIN rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 455.630 0.460 456.090 ;
    END
  END rd_out[290]
  PIN rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 456.090 0.460 456.550 ;
    END
  END rd_out[291]
  PIN rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 456.550 0.460 457.010 ;
    END
  END rd_out[292]
  PIN rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 457.010 0.460 457.470 ;
    END
  END rd_out[293]
  PIN rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 457.470 0.460 457.930 ;
    END
  END rd_out[294]
  PIN rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 457.930 0.460 458.390 ;
    END
  END rd_out[295]
  PIN rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 458.390 0.460 458.850 ;
    END
  END rd_out[296]
  PIN rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 458.850 0.460 459.310 ;
    END
  END rd_out[297]
  PIN rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 459.310 0.460 459.770 ;
    END
  END rd_out[298]
  PIN rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 459.770 0.460 460.230 ;
    END
  END rd_out[299]
  PIN rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 460.230 0.460 460.690 ;
    END
  END rd_out[300]
  PIN rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 460.690 0.460 461.150 ;
    END
  END rd_out[301]
  PIN rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 461.150 0.460 461.610 ;
    END
  END rd_out[302]
  PIN rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 461.610 0.460 462.070 ;
    END
  END rd_out[303]
  PIN rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 462.070 0.460 462.530 ;
    END
  END rd_out[304]
  PIN rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 462.530 0.460 462.990 ;
    END
  END rd_out[305]
  PIN rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 462.990 0.460 463.450 ;
    END
  END rd_out[306]
  PIN rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 463.450 0.460 463.910 ;
    END
  END rd_out[307]
  PIN rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 463.910 0.460 464.370 ;
    END
  END rd_out[308]
  PIN rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 464.370 0.460 464.830 ;
    END
  END rd_out[309]
  PIN rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 464.830 0.460 465.290 ;
    END
  END rd_out[310]
  PIN rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 465.290 0.460 465.750 ;
    END
  END rd_out[311]
  PIN rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 465.750 0.460 466.210 ;
    END
  END rd_out[312]
  PIN rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 466.210 0.460 466.670 ;
    END
  END rd_out[313]
  PIN rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 466.670 0.460 467.130 ;
    END
  END rd_out[314]
  PIN rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 467.130 0.460 467.590 ;
    END
  END rd_out[315]
  PIN rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 467.590 0.460 468.050 ;
    END
  END rd_out[316]
  PIN rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 468.050 0.460 468.510 ;
    END
  END rd_out[317]
  PIN rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 468.510 0.460 468.970 ;
    END
  END rd_out[318]
  PIN rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 468.970 0.460 469.430 ;
    END
  END rd_out[319]
  PIN rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 469.430 0.460 469.890 ;
    END
  END rd_out[320]
  PIN rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 469.890 0.460 470.350 ;
    END
  END rd_out[321]
  PIN rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 470.350 0.460 470.810 ;
    END
  END rd_out[322]
  PIN rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 470.810 0.460 471.270 ;
    END
  END rd_out[323]
  PIN rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 471.270 0.460 471.730 ;
    END
  END rd_out[324]
  PIN rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 471.730 0.460 472.190 ;
    END
  END rd_out[325]
  PIN rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 472.190 0.460 472.650 ;
    END
  END rd_out[326]
  PIN rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 472.650 0.460 473.110 ;
    END
  END rd_out[327]
  PIN rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 473.110 0.460 473.570 ;
    END
  END rd_out[328]
  PIN rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 473.570 0.460 474.030 ;
    END
  END rd_out[329]
  PIN rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 474.030 0.460 474.490 ;
    END
  END rd_out[330]
  PIN rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 474.490 0.460 474.950 ;
    END
  END rd_out[331]
  PIN rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 474.950 0.460 475.410 ;
    END
  END rd_out[332]
  PIN rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 475.410 0.460 475.870 ;
    END
  END rd_out[333]
  PIN rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 475.870 0.460 476.330 ;
    END
  END rd_out[334]
  PIN rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 476.330 0.460 476.790 ;
    END
  END rd_out[335]
  PIN rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 476.790 0.460 477.250 ;
    END
  END rd_out[336]
  PIN rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 477.250 0.460 477.710 ;
    END
  END rd_out[337]
  PIN rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 477.710 0.460 478.170 ;
    END
  END rd_out[338]
  PIN rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 478.170 0.460 478.630 ;
    END
  END rd_out[339]
  PIN rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 478.630 0.460 479.090 ;
    END
  END rd_out[340]
  PIN rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 479.090 0.460 479.550 ;
    END
  END rd_out[341]
  PIN rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 479.550 0.460 480.010 ;
    END
  END rd_out[342]
  PIN rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 480.010 0.460 480.470 ;
    END
  END rd_out[343]
  PIN rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 480.470 0.460 480.930 ;
    END
  END rd_out[344]
  PIN rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 480.930 0.460 481.390 ;
    END
  END rd_out[345]
  PIN rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 481.390 0.460 481.850 ;
    END
  END rd_out[346]
  PIN rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 481.850 0.460 482.310 ;
    END
  END rd_out[347]
  PIN rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 482.310 0.460 482.770 ;
    END
  END rd_out[348]
  PIN rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 482.770 0.460 483.230 ;
    END
  END rd_out[349]
  PIN rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 483.230 0.460 483.690 ;
    END
  END rd_out[350]
  PIN rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 483.690 0.460 484.150 ;
    END
  END rd_out[351]
  PIN rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 484.150 0.460 484.610 ;
    END
  END rd_out[352]
  PIN rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 484.610 0.460 485.070 ;
    END
  END rd_out[353]
  PIN rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.070 0.460 485.530 ;
    END
  END rd_out[354]
  PIN rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.530 0.460 485.990 ;
    END
  END rd_out[355]
  PIN rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.990 0.460 486.450 ;
    END
  END rd_out[356]
  PIN rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 486.450 0.460 486.910 ;
    END
  END rd_out[357]
  PIN rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 486.910 0.460 487.370 ;
    END
  END rd_out[358]
  PIN rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 487.370 0.460 487.830 ;
    END
  END rd_out[359]
  PIN rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 487.830 0.460 488.290 ;
    END
  END rd_out[360]
  PIN rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 488.290 0.460 488.750 ;
    END
  END rd_out[361]
  PIN rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 488.750 0.460 489.210 ;
    END
  END rd_out[362]
  PIN rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 489.210 0.460 489.670 ;
    END
  END rd_out[363]
  PIN rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 489.670 0.460 490.130 ;
    END
  END rd_out[364]
  PIN rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 490.130 0.460 490.590 ;
    END
  END rd_out[365]
  PIN rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 490.590 0.460 491.050 ;
    END
  END rd_out[366]
  PIN rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 491.050 0.460 491.510 ;
    END
  END rd_out[367]
  PIN rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 491.510 0.460 491.970 ;
    END
  END rd_out[368]
  PIN rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 491.970 0.460 492.430 ;
    END
  END rd_out[369]
  PIN rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 492.430 0.460 492.890 ;
    END
  END rd_out[370]
  PIN rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 492.890 0.460 493.350 ;
    END
  END rd_out[371]
  PIN rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 493.350 0.460 493.810 ;
    END
  END rd_out[372]
  PIN rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 493.810 0.460 494.270 ;
    END
  END rd_out[373]
  PIN rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 494.270 0.460 494.730 ;
    END
  END rd_out[374]
  PIN rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 494.730 0.460 495.190 ;
    END
  END rd_out[375]
  PIN rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 495.190 0.460 495.650 ;
    END
  END rd_out[376]
  PIN rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 495.650 0.460 496.110 ;
    END
  END rd_out[377]
  PIN rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 496.110 0.460 496.570 ;
    END
  END rd_out[378]
  PIN rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 496.570 0.460 497.030 ;
    END
  END rd_out[379]
  PIN rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 497.030 0.460 497.490 ;
    END
  END rd_out[380]
  PIN rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 497.490 0.460 497.950 ;
    END
  END rd_out[381]
  PIN rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 497.950 0.460 498.410 ;
    END
  END rd_out[382]
  PIN rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 498.410 0.460 498.870 ;
    END
  END rd_out[383]
  PIN rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 498.870 0.460 499.330 ;
    END
  END rd_out[384]
  PIN rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 499.330 0.460 499.790 ;
    END
  END rd_out[385]
  PIN rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 499.790 0.460 500.250 ;
    END
  END rd_out[386]
  PIN rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 500.250 0.460 500.710 ;
    END
  END rd_out[387]
  PIN rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 500.710 0.460 501.170 ;
    END
  END rd_out[388]
  PIN rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.170 0.460 501.630 ;
    END
  END rd_out[389]
  PIN rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.630 0.460 502.090 ;
    END
  END rd_out[390]
  PIN rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 502.090 0.460 502.550 ;
    END
  END rd_out[391]
  PIN rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 502.550 0.460 503.010 ;
    END
  END rd_out[392]
  PIN rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 503.010 0.460 503.470 ;
    END
  END rd_out[393]
  PIN rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 503.470 0.460 503.930 ;
    END
  END rd_out[394]
  PIN rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 503.930 0.460 504.390 ;
    END
  END rd_out[395]
  PIN rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 504.390 0.460 504.850 ;
    END
  END rd_out[396]
  PIN rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 504.850 0.460 505.310 ;
    END
  END rd_out[397]
  PIN rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 505.310 0.460 505.770 ;
    END
  END rd_out[398]
  PIN rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 505.770 0.460 506.230 ;
    END
  END rd_out[399]
  PIN rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 506.230 0.460 506.690 ;
    END
  END rd_out[400]
  PIN rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 506.690 0.460 507.150 ;
    END
  END rd_out[401]
  PIN rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 507.150 0.460 507.610 ;
    END
  END rd_out[402]
  PIN rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 507.610 0.460 508.070 ;
    END
  END rd_out[403]
  PIN rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 508.070 0.460 508.530 ;
    END
  END rd_out[404]
  PIN rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 508.530 0.460 508.990 ;
    END
  END rd_out[405]
  PIN rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 508.990 0.460 509.450 ;
    END
  END rd_out[406]
  PIN rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 509.450 0.460 509.910 ;
    END
  END rd_out[407]
  PIN rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 509.910 0.460 510.370 ;
    END
  END rd_out[408]
  PIN rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 510.370 0.460 510.830 ;
    END
  END rd_out[409]
  PIN rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 510.830 0.460 511.290 ;
    END
  END rd_out[410]
  PIN rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 511.290 0.460 511.750 ;
    END
  END rd_out[411]
  PIN rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 511.750 0.460 512.210 ;
    END
  END rd_out[412]
  PIN rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 512.210 0.460 512.670 ;
    END
  END rd_out[413]
  PIN rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 512.670 0.460 513.130 ;
    END
  END rd_out[414]
  PIN rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 513.130 0.460 513.590 ;
    END
  END rd_out[415]
  PIN rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 513.590 0.460 514.050 ;
    END
  END rd_out[416]
  PIN rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 514.050 0.460 514.510 ;
    END
  END rd_out[417]
  PIN rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 514.510 0.460 514.970 ;
    END
  END rd_out[418]
  PIN rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 514.970 0.460 515.430 ;
    END
  END rd_out[419]
  PIN rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 515.430 0.460 515.890 ;
    END
  END rd_out[420]
  PIN rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 515.890 0.460 516.350 ;
    END
  END rd_out[421]
  PIN rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 516.350 0.460 516.810 ;
    END
  END rd_out[422]
  PIN rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 516.810 0.460 517.270 ;
    END
  END rd_out[423]
  PIN rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 517.270 0.460 517.730 ;
    END
  END rd_out[424]
  PIN rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 517.730 0.460 518.190 ;
    END
  END rd_out[425]
  PIN rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 518.190 0.460 518.650 ;
    END
  END rd_out[426]
  PIN rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 518.650 0.460 519.110 ;
    END
  END rd_out[427]
  PIN rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 519.110 0.460 519.570 ;
    END
  END rd_out[428]
  PIN rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 519.570 0.460 520.030 ;
    END
  END rd_out[429]
  PIN rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 520.030 0.460 520.490 ;
    END
  END rd_out[430]
  PIN rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 520.490 0.460 520.950 ;
    END
  END rd_out[431]
  PIN rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 520.950 0.460 521.410 ;
    END
  END rd_out[432]
  PIN rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 521.410 0.460 521.870 ;
    END
  END rd_out[433]
  PIN rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 521.870 0.460 522.330 ;
    END
  END rd_out[434]
  PIN rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 522.330 0.460 522.790 ;
    END
  END rd_out[435]
  PIN rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 522.790 0.460 523.250 ;
    END
  END rd_out[436]
  PIN rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 523.250 0.460 523.710 ;
    END
  END rd_out[437]
  PIN rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 523.710 0.460 524.170 ;
    END
  END rd_out[438]
  PIN rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 524.170 0.460 524.630 ;
    END
  END rd_out[439]
  PIN rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 524.630 0.460 525.090 ;
    END
  END rd_out[440]
  PIN rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 525.090 0.460 525.550 ;
    END
  END rd_out[441]
  PIN rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 525.550 0.460 526.010 ;
    END
  END rd_out[442]
  PIN rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.010 0.460 526.470 ;
    END
  END rd_out[443]
  PIN rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.470 0.460 526.930 ;
    END
  END rd_out[444]
  PIN rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.930 0.460 527.390 ;
    END
  END rd_out[445]
  PIN rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 527.390 0.460 527.850 ;
    END
  END rd_out[446]
  PIN rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 527.850 0.460 528.310 ;
    END
  END rd_out[447]
  PIN rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 528.310 0.460 528.770 ;
    END
  END rd_out[448]
  PIN rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 528.770 0.460 529.230 ;
    END
  END rd_out[449]
  PIN rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 529.230 0.460 529.690 ;
    END
  END rd_out[450]
  PIN rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 529.690 0.460 530.150 ;
    END
  END rd_out[451]
  PIN rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 530.150 0.460 530.610 ;
    END
  END rd_out[452]
  PIN rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 530.610 0.460 531.070 ;
    END
  END rd_out[453]
  PIN rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 531.070 0.460 531.530 ;
    END
  END rd_out[454]
  PIN rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 531.530 0.460 531.990 ;
    END
  END rd_out[455]
  PIN rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 531.990 0.460 532.450 ;
    END
  END rd_out[456]
  PIN rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 532.450 0.460 532.910 ;
    END
  END rd_out[457]
  PIN rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 532.910 0.460 533.370 ;
    END
  END rd_out[458]
  PIN rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 533.370 0.460 533.830 ;
    END
  END rd_out[459]
  PIN rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 533.830 0.460 534.290 ;
    END
  END rd_out[460]
  PIN rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 534.290 0.460 534.750 ;
    END
  END rd_out[461]
  PIN rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 534.750 0.460 535.210 ;
    END
  END rd_out[462]
  PIN rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.210 0.460 535.670 ;
    END
  END rd_out[463]
  PIN rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.670 0.460 536.130 ;
    END
  END rd_out[464]
  PIN rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 536.130 0.460 536.590 ;
    END
  END rd_out[465]
  PIN rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 536.590 0.460 537.050 ;
    END
  END rd_out[466]
  PIN rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 537.050 0.460 537.510 ;
    END
  END rd_out[467]
  PIN rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 537.510 0.460 537.970 ;
    END
  END rd_out[468]
  PIN rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 537.970 0.460 538.430 ;
    END
  END rd_out[469]
  PIN rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 538.430 0.460 538.890 ;
    END
  END rd_out[470]
  PIN rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 538.890 0.460 539.350 ;
    END
  END rd_out[471]
  PIN rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 539.350 0.460 539.810 ;
    END
  END rd_out[472]
  PIN rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 539.810 0.460 540.270 ;
    END
  END rd_out[473]
  PIN rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 540.270 0.460 540.730 ;
    END
  END rd_out[474]
  PIN rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 540.730 0.460 541.190 ;
    END
  END rd_out[475]
  PIN rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 541.190 0.460 541.650 ;
    END
  END rd_out[476]
  PIN rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 541.650 0.460 542.110 ;
    END
  END rd_out[477]
  PIN rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 542.110 0.460 542.570 ;
    END
  END rd_out[478]
  PIN rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 542.570 0.460 543.030 ;
    END
  END rd_out[479]
  PIN rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.030 0.460 543.490 ;
    END
  END rd_out[480]
  PIN rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.490 0.460 543.950 ;
    END
  END rd_out[481]
  PIN rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.950 0.460 544.410 ;
    END
  END rd_out[482]
  PIN rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 544.410 0.460 544.870 ;
    END
  END rd_out[483]
  PIN rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 544.870 0.460 545.330 ;
    END
  END rd_out[484]
  PIN rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 545.330 0.460 545.790 ;
    END
  END rd_out[485]
  PIN rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 545.790 0.460 546.250 ;
    END
  END rd_out[486]
  PIN rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 546.250 0.460 546.710 ;
    END
  END rd_out[487]
  PIN rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 546.710 0.460 547.170 ;
    END
  END rd_out[488]
  PIN rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 547.170 0.460 547.630 ;
    END
  END rd_out[489]
  PIN rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 547.630 0.460 548.090 ;
    END
  END rd_out[490]
  PIN rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 548.090 0.460 548.550 ;
    END
  END rd_out[491]
  PIN rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 548.550 0.460 549.010 ;
    END
  END rd_out[492]
  PIN rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 549.010 0.460 549.470 ;
    END
  END rd_out[493]
  PIN rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 549.470 0.460 549.930 ;
    END
  END rd_out[494]
  PIN rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 549.930 0.460 550.390 ;
    END
  END rd_out[495]
  PIN rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 550.390 0.460 550.850 ;
    END
  END rd_out[496]
  PIN rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 550.850 0.460 551.310 ;
    END
  END rd_out[497]
  PIN rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 551.310 0.460 551.770 ;
    END
  END rd_out[498]
  PIN rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 551.770 0.460 552.230 ;
    END
  END rd_out[499]
  PIN rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 552.230 0.460 552.690 ;
    END
  END rd_out[500]
  PIN rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 552.690 0.460 553.150 ;
    END
  END rd_out[501]
  PIN rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 553.150 0.460 553.610 ;
    END
  END rd_out[502]
  PIN rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 553.610 0.460 554.070 ;
    END
  END rd_out[503]
  PIN rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 554.070 0.460 554.530 ;
    END
  END rd_out[504]
  PIN rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 554.530 0.460 554.990 ;
    END
  END rd_out[505]
  PIN rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 554.990 0.460 555.450 ;
    END
  END rd_out[506]
  PIN rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 555.450 0.460 555.910 ;
    END
  END rd_out[507]
  PIN rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 555.910 0.460 556.370 ;
    END
  END rd_out[508]
  PIN rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 556.370 0.460 556.830 ;
    END
  END rd_out[509]
  PIN rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 556.830 0.460 557.290 ;
    END
  END rd_out[510]
  PIN rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 557.290 0.460 557.750 ;
    END
  END rd_out[511]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 640.090 0.460 640.550 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 640.550 0.460 641.010 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 641.010 0.460 641.470 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 641.470 0.460 641.930 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 641.930 0.460 642.390 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 642.390 0.460 642.850 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 642.850 0.460 643.310 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 643.310 0.460 643.770 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 643.770 0.460 644.230 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 644.230 0.460 644.690 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 644.690 0.460 645.150 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 645.150 0.460 645.610 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 645.610 0.460 646.070 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 646.070 0.460 646.530 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 646.530 0.460 646.990 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 646.990 0.460 647.450 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 647.450 0.460 647.910 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 647.910 0.460 648.370 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 648.370 0.460 648.830 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 648.830 0.460 649.290 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 649.290 0.460 649.750 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 649.750 0.460 650.210 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 650.210 0.460 650.670 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 650.670 0.460 651.130 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 651.130 0.460 651.590 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 651.590 0.460 652.050 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 652.050 0.460 652.510 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 652.510 0.460 652.970 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 652.970 0.460 653.430 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 653.430 0.460 653.890 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 653.890 0.460 654.350 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 654.350 0.460 654.810 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 654.810 0.460 655.270 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 655.270 0.460 655.730 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 655.730 0.460 656.190 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 656.190 0.460 656.650 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 656.650 0.460 657.110 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 657.110 0.460 657.570 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 657.570 0.460 658.030 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 658.030 0.460 658.490 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 658.490 0.460 658.950 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 658.950 0.460 659.410 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 659.410 0.460 659.870 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 659.870 0.460 660.330 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 660.330 0.460 660.790 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 660.790 0.460 661.250 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 661.250 0.460 661.710 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 661.710 0.460 662.170 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 662.170 0.460 662.630 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 662.630 0.460 663.090 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 663.090 0.460 663.550 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 663.550 0.460 664.010 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 664.010 0.460 664.470 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 664.470 0.460 664.930 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 664.930 0.460 665.390 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 665.390 0.460 665.850 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 665.850 0.460 666.310 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 666.310 0.460 666.770 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 666.770 0.460 667.230 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 667.230 0.460 667.690 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 667.690 0.460 668.150 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 668.150 0.460 668.610 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 668.610 0.460 669.070 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 669.070 0.460 669.530 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 669.530 0.460 669.990 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 669.990 0.460 670.450 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 670.450 0.460 670.910 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 670.910 0.460 671.370 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 671.370 0.460 671.830 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 671.830 0.460 672.290 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 672.290 0.460 672.750 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 672.750 0.460 673.210 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 673.210 0.460 673.670 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 673.670 0.460 674.130 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 674.130 0.460 674.590 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 674.590 0.460 675.050 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 675.050 0.460 675.510 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 675.510 0.460 675.970 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 675.970 0.460 676.430 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 676.430 0.460 676.890 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 676.890 0.460 677.350 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 677.350 0.460 677.810 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 677.810 0.460 678.270 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 678.270 0.460 678.730 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 678.730 0.460 679.190 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 679.190 0.460 679.650 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 679.650 0.460 680.110 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 680.110 0.460 680.570 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 680.570 0.460 681.030 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 681.030 0.460 681.490 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 681.490 0.460 681.950 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 681.950 0.460 682.410 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 682.410 0.460 682.870 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 682.870 0.460 683.330 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 683.330 0.460 683.790 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 683.790 0.460 684.250 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 684.250 0.460 684.710 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 684.710 0.460 685.170 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 685.170 0.460 685.630 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 685.630 0.460 686.090 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 686.090 0.460 686.550 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 686.550 0.460 687.010 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 687.010 0.460 687.470 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 687.470 0.460 687.930 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 687.930 0.460 688.390 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 688.390 0.460 688.850 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 688.850 0.460 689.310 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 689.310 0.460 689.770 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 689.770 0.460 690.230 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 690.230 0.460 690.690 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 690.690 0.460 691.150 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 691.150 0.460 691.610 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 691.610 0.460 692.070 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 692.070 0.460 692.530 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 692.530 0.460 692.990 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 692.990 0.460 693.450 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 693.450 0.460 693.910 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 693.910 0.460 694.370 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 694.370 0.460 694.830 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 694.830 0.460 695.290 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 695.290 0.460 695.750 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 695.750 0.460 696.210 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 696.210 0.460 696.670 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 696.670 0.460 697.130 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 697.130 0.460 697.590 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 697.590 0.460 698.050 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 698.050 0.460 698.510 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 698.510 0.460 698.970 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 698.970 0.460 699.430 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 699.430 0.460 699.890 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 699.890 0.460 700.350 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 700.350 0.460 700.810 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 700.810 0.460 701.270 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 701.270 0.460 701.730 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 701.730 0.460 702.190 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 702.190 0.460 702.650 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 702.650 0.460 703.110 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 703.110 0.460 703.570 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 703.570 0.460 704.030 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 704.030 0.460 704.490 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 704.490 0.460 704.950 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 704.950 0.460 705.410 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 705.410 0.460 705.870 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 705.870 0.460 706.330 ;
    END
  END wd_in[143]
  PIN wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 706.330 0.460 706.790 ;
    END
  END wd_in[144]
  PIN wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 706.790 0.460 707.250 ;
    END
  END wd_in[145]
  PIN wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 707.250 0.460 707.710 ;
    END
  END wd_in[146]
  PIN wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 707.710 0.460 708.170 ;
    END
  END wd_in[147]
  PIN wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 708.170 0.460 708.630 ;
    END
  END wd_in[148]
  PIN wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 708.630 0.460 709.090 ;
    END
  END wd_in[149]
  PIN wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 709.090 0.460 709.550 ;
    END
  END wd_in[150]
  PIN wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 709.550 0.460 710.010 ;
    END
  END wd_in[151]
  PIN wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 710.010 0.460 710.470 ;
    END
  END wd_in[152]
  PIN wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 710.470 0.460 710.930 ;
    END
  END wd_in[153]
  PIN wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 710.930 0.460 711.390 ;
    END
  END wd_in[154]
  PIN wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 711.390 0.460 711.850 ;
    END
  END wd_in[155]
  PIN wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 711.850 0.460 712.310 ;
    END
  END wd_in[156]
  PIN wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 712.310 0.460 712.770 ;
    END
  END wd_in[157]
  PIN wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 712.770 0.460 713.230 ;
    END
  END wd_in[158]
  PIN wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 713.230 0.460 713.690 ;
    END
  END wd_in[159]
  PIN wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 713.690 0.460 714.150 ;
    END
  END wd_in[160]
  PIN wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 714.150 0.460 714.610 ;
    END
  END wd_in[161]
  PIN wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 714.610 0.460 715.070 ;
    END
  END wd_in[162]
  PIN wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 715.070 0.460 715.530 ;
    END
  END wd_in[163]
  PIN wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 715.530 0.460 715.990 ;
    END
  END wd_in[164]
  PIN wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 715.990 0.460 716.450 ;
    END
  END wd_in[165]
  PIN wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 716.450 0.460 716.910 ;
    END
  END wd_in[166]
  PIN wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 716.910 0.460 717.370 ;
    END
  END wd_in[167]
  PIN wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 717.370 0.460 717.830 ;
    END
  END wd_in[168]
  PIN wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 717.830 0.460 718.290 ;
    END
  END wd_in[169]
  PIN wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 718.290 0.460 718.750 ;
    END
  END wd_in[170]
  PIN wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 718.750 0.460 719.210 ;
    END
  END wd_in[171]
  PIN wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 719.210 0.460 719.670 ;
    END
  END wd_in[172]
  PIN wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 719.670 0.460 720.130 ;
    END
  END wd_in[173]
  PIN wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 720.130 0.460 720.590 ;
    END
  END wd_in[174]
  PIN wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 720.590 0.460 721.050 ;
    END
  END wd_in[175]
  PIN wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 721.050 0.460 721.510 ;
    END
  END wd_in[176]
  PIN wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 721.510 0.460 721.970 ;
    END
  END wd_in[177]
  PIN wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 721.970 0.460 722.430 ;
    END
  END wd_in[178]
  PIN wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 722.430 0.460 722.890 ;
    END
  END wd_in[179]
  PIN wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 722.890 0.460 723.350 ;
    END
  END wd_in[180]
  PIN wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 723.350 0.460 723.810 ;
    END
  END wd_in[181]
  PIN wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 723.810 0.460 724.270 ;
    END
  END wd_in[182]
  PIN wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 724.270 0.460 724.730 ;
    END
  END wd_in[183]
  PIN wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 724.730 0.460 725.190 ;
    END
  END wd_in[184]
  PIN wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 725.190 0.460 725.650 ;
    END
  END wd_in[185]
  PIN wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 725.650 0.460 726.110 ;
    END
  END wd_in[186]
  PIN wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 726.110 0.460 726.570 ;
    END
  END wd_in[187]
  PIN wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 726.570 0.460 727.030 ;
    END
  END wd_in[188]
  PIN wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 727.030 0.460 727.490 ;
    END
  END wd_in[189]
  PIN wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 727.490 0.460 727.950 ;
    END
  END wd_in[190]
  PIN wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 727.950 0.460 728.410 ;
    END
  END wd_in[191]
  PIN wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 728.410 0.460 728.870 ;
    END
  END wd_in[192]
  PIN wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 728.870 0.460 729.330 ;
    END
  END wd_in[193]
  PIN wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 729.330 0.460 729.790 ;
    END
  END wd_in[194]
  PIN wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 729.790 0.460 730.250 ;
    END
  END wd_in[195]
  PIN wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 730.250 0.460 730.710 ;
    END
  END wd_in[196]
  PIN wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 730.710 0.460 731.170 ;
    END
  END wd_in[197]
  PIN wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 731.170 0.460 731.630 ;
    END
  END wd_in[198]
  PIN wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 731.630 0.460 732.090 ;
    END
  END wd_in[199]
  PIN wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 732.090 0.460 732.550 ;
    END
  END wd_in[200]
  PIN wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 732.550 0.460 733.010 ;
    END
  END wd_in[201]
  PIN wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 733.010 0.460 733.470 ;
    END
  END wd_in[202]
  PIN wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 733.470 0.460 733.930 ;
    END
  END wd_in[203]
  PIN wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 733.930 0.460 734.390 ;
    END
  END wd_in[204]
  PIN wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 734.390 0.460 734.850 ;
    END
  END wd_in[205]
  PIN wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 734.850 0.460 735.310 ;
    END
  END wd_in[206]
  PIN wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 735.310 0.460 735.770 ;
    END
  END wd_in[207]
  PIN wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 735.770 0.460 736.230 ;
    END
  END wd_in[208]
  PIN wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 736.230 0.460 736.690 ;
    END
  END wd_in[209]
  PIN wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 736.690 0.460 737.150 ;
    END
  END wd_in[210]
  PIN wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 737.150 0.460 737.610 ;
    END
  END wd_in[211]
  PIN wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 737.610 0.460 738.070 ;
    END
  END wd_in[212]
  PIN wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 738.070 0.460 738.530 ;
    END
  END wd_in[213]
  PIN wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 738.530 0.460 738.990 ;
    END
  END wd_in[214]
  PIN wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 738.990 0.460 739.450 ;
    END
  END wd_in[215]
  PIN wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 739.450 0.460 739.910 ;
    END
  END wd_in[216]
  PIN wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 739.910 0.460 740.370 ;
    END
  END wd_in[217]
  PIN wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 740.370 0.460 740.830 ;
    END
  END wd_in[218]
  PIN wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 740.830 0.460 741.290 ;
    END
  END wd_in[219]
  PIN wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 741.290 0.460 741.750 ;
    END
  END wd_in[220]
  PIN wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 741.750 0.460 742.210 ;
    END
  END wd_in[221]
  PIN wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 742.210 0.460 742.670 ;
    END
  END wd_in[222]
  PIN wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 742.670 0.460 743.130 ;
    END
  END wd_in[223]
  PIN wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 743.130 0.460 743.590 ;
    END
  END wd_in[224]
  PIN wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 743.590 0.460 744.050 ;
    END
  END wd_in[225]
  PIN wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 744.050 0.460 744.510 ;
    END
  END wd_in[226]
  PIN wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 744.510 0.460 744.970 ;
    END
  END wd_in[227]
  PIN wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 744.970 0.460 745.430 ;
    END
  END wd_in[228]
  PIN wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 745.430 0.460 745.890 ;
    END
  END wd_in[229]
  PIN wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 745.890 0.460 746.350 ;
    END
  END wd_in[230]
  PIN wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 746.350 0.460 746.810 ;
    END
  END wd_in[231]
  PIN wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 746.810 0.460 747.270 ;
    END
  END wd_in[232]
  PIN wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 747.270 0.460 747.730 ;
    END
  END wd_in[233]
  PIN wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 747.730 0.460 748.190 ;
    END
  END wd_in[234]
  PIN wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 748.190 0.460 748.650 ;
    END
  END wd_in[235]
  PIN wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 748.650 0.460 749.110 ;
    END
  END wd_in[236]
  PIN wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 749.110 0.460 749.570 ;
    END
  END wd_in[237]
  PIN wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 749.570 0.460 750.030 ;
    END
  END wd_in[238]
  PIN wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 750.030 0.460 750.490 ;
    END
  END wd_in[239]
  PIN wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 750.490 0.460 750.950 ;
    END
  END wd_in[240]
  PIN wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 750.950 0.460 751.410 ;
    END
  END wd_in[241]
  PIN wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 751.410 0.460 751.870 ;
    END
  END wd_in[242]
  PIN wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 751.870 0.460 752.330 ;
    END
  END wd_in[243]
  PIN wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 752.330 0.460 752.790 ;
    END
  END wd_in[244]
  PIN wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 752.790 0.460 753.250 ;
    END
  END wd_in[245]
  PIN wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 753.250 0.460 753.710 ;
    END
  END wd_in[246]
  PIN wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 753.710 0.460 754.170 ;
    END
  END wd_in[247]
  PIN wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 754.170 0.460 754.630 ;
    END
  END wd_in[248]
  PIN wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 754.630 0.460 755.090 ;
    END
  END wd_in[249]
  PIN wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 755.090 0.460 755.550 ;
    END
  END wd_in[250]
  PIN wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 755.550 0.460 756.010 ;
    END
  END wd_in[251]
  PIN wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 756.010 0.460 756.470 ;
    END
  END wd_in[252]
  PIN wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 756.470 0.460 756.930 ;
    END
  END wd_in[253]
  PIN wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 756.930 0.460 757.390 ;
    END
  END wd_in[254]
  PIN wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 757.390 0.460 757.850 ;
    END
  END wd_in[255]
  PIN wd_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 757.850 0.460 758.310 ;
    END
  END wd_in[256]
  PIN wd_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 758.310 0.460 758.770 ;
    END
  END wd_in[257]
  PIN wd_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 758.770 0.460 759.230 ;
    END
  END wd_in[258]
  PIN wd_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 759.230 0.460 759.690 ;
    END
  END wd_in[259]
  PIN wd_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 759.690 0.460 760.150 ;
    END
  END wd_in[260]
  PIN wd_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 760.150 0.460 760.610 ;
    END
  END wd_in[261]
  PIN wd_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 760.610 0.460 761.070 ;
    END
  END wd_in[262]
  PIN wd_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 761.070 0.460 761.530 ;
    END
  END wd_in[263]
  PIN wd_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 761.530 0.460 761.990 ;
    END
  END wd_in[264]
  PIN wd_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 761.990 0.460 762.450 ;
    END
  END wd_in[265]
  PIN wd_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 762.450 0.460 762.910 ;
    END
  END wd_in[266]
  PIN wd_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 762.910 0.460 763.370 ;
    END
  END wd_in[267]
  PIN wd_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 763.370 0.460 763.830 ;
    END
  END wd_in[268]
  PIN wd_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 763.830 0.460 764.290 ;
    END
  END wd_in[269]
  PIN wd_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 764.290 0.460 764.750 ;
    END
  END wd_in[270]
  PIN wd_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 764.750 0.460 765.210 ;
    END
  END wd_in[271]
  PIN wd_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 765.210 0.460 765.670 ;
    END
  END wd_in[272]
  PIN wd_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 765.670 0.460 766.130 ;
    END
  END wd_in[273]
  PIN wd_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 766.130 0.460 766.590 ;
    END
  END wd_in[274]
  PIN wd_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 766.590 0.460 767.050 ;
    END
  END wd_in[275]
  PIN wd_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 767.050 0.460 767.510 ;
    END
  END wd_in[276]
  PIN wd_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 767.510 0.460 767.970 ;
    END
  END wd_in[277]
  PIN wd_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 767.970 0.460 768.430 ;
    END
  END wd_in[278]
  PIN wd_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 768.430 0.460 768.890 ;
    END
  END wd_in[279]
  PIN wd_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 768.890 0.460 769.350 ;
    END
  END wd_in[280]
  PIN wd_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 769.350 0.460 769.810 ;
    END
  END wd_in[281]
  PIN wd_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 769.810 0.460 770.270 ;
    END
  END wd_in[282]
  PIN wd_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 770.270 0.460 770.730 ;
    END
  END wd_in[283]
  PIN wd_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 770.730 0.460 771.190 ;
    END
  END wd_in[284]
  PIN wd_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 771.190 0.460 771.650 ;
    END
  END wd_in[285]
  PIN wd_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 771.650 0.460 772.110 ;
    END
  END wd_in[286]
  PIN wd_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 772.110 0.460 772.570 ;
    END
  END wd_in[287]
  PIN wd_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 772.570 0.460 773.030 ;
    END
  END wd_in[288]
  PIN wd_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 773.030 0.460 773.490 ;
    END
  END wd_in[289]
  PIN wd_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 773.490 0.460 773.950 ;
    END
  END wd_in[290]
  PIN wd_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 773.950 0.460 774.410 ;
    END
  END wd_in[291]
  PIN wd_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 774.410 0.460 774.870 ;
    END
  END wd_in[292]
  PIN wd_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 774.870 0.460 775.330 ;
    END
  END wd_in[293]
  PIN wd_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 775.330 0.460 775.790 ;
    END
  END wd_in[294]
  PIN wd_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 775.790 0.460 776.250 ;
    END
  END wd_in[295]
  PIN wd_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 776.250 0.460 776.710 ;
    END
  END wd_in[296]
  PIN wd_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 776.710 0.460 777.170 ;
    END
  END wd_in[297]
  PIN wd_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 777.170 0.460 777.630 ;
    END
  END wd_in[298]
  PIN wd_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 777.630 0.460 778.090 ;
    END
  END wd_in[299]
  PIN wd_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 778.090 0.460 778.550 ;
    END
  END wd_in[300]
  PIN wd_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 778.550 0.460 779.010 ;
    END
  END wd_in[301]
  PIN wd_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 779.010 0.460 779.470 ;
    END
  END wd_in[302]
  PIN wd_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 779.470 0.460 779.930 ;
    END
  END wd_in[303]
  PIN wd_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 779.930 0.460 780.390 ;
    END
  END wd_in[304]
  PIN wd_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 780.390 0.460 780.850 ;
    END
  END wd_in[305]
  PIN wd_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 780.850 0.460 781.310 ;
    END
  END wd_in[306]
  PIN wd_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 781.310 0.460 781.770 ;
    END
  END wd_in[307]
  PIN wd_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 781.770 0.460 782.230 ;
    END
  END wd_in[308]
  PIN wd_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 782.230 0.460 782.690 ;
    END
  END wd_in[309]
  PIN wd_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 782.690 0.460 783.150 ;
    END
  END wd_in[310]
  PIN wd_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 783.150 0.460 783.610 ;
    END
  END wd_in[311]
  PIN wd_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 783.610 0.460 784.070 ;
    END
  END wd_in[312]
  PIN wd_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 784.070 0.460 784.530 ;
    END
  END wd_in[313]
  PIN wd_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 784.530 0.460 784.990 ;
    END
  END wd_in[314]
  PIN wd_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 784.990 0.460 785.450 ;
    END
  END wd_in[315]
  PIN wd_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 785.450 0.460 785.910 ;
    END
  END wd_in[316]
  PIN wd_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 785.910 0.460 786.370 ;
    END
  END wd_in[317]
  PIN wd_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 786.370 0.460 786.830 ;
    END
  END wd_in[318]
  PIN wd_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 786.830 0.460 787.290 ;
    END
  END wd_in[319]
  PIN wd_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 787.290 0.460 787.750 ;
    END
  END wd_in[320]
  PIN wd_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 787.750 0.460 788.210 ;
    END
  END wd_in[321]
  PIN wd_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 788.210 0.460 788.670 ;
    END
  END wd_in[322]
  PIN wd_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 788.670 0.460 789.130 ;
    END
  END wd_in[323]
  PIN wd_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 789.130 0.460 789.590 ;
    END
  END wd_in[324]
  PIN wd_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 789.590 0.460 790.050 ;
    END
  END wd_in[325]
  PIN wd_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 790.050 0.460 790.510 ;
    END
  END wd_in[326]
  PIN wd_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 790.510 0.460 790.970 ;
    END
  END wd_in[327]
  PIN wd_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 790.970 0.460 791.430 ;
    END
  END wd_in[328]
  PIN wd_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 791.430 0.460 791.890 ;
    END
  END wd_in[329]
  PIN wd_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 791.890 0.460 792.350 ;
    END
  END wd_in[330]
  PIN wd_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 792.350 0.460 792.810 ;
    END
  END wd_in[331]
  PIN wd_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 792.810 0.460 793.270 ;
    END
  END wd_in[332]
  PIN wd_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 793.270 0.460 793.730 ;
    END
  END wd_in[333]
  PIN wd_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 793.730 0.460 794.190 ;
    END
  END wd_in[334]
  PIN wd_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 794.190 0.460 794.650 ;
    END
  END wd_in[335]
  PIN wd_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 794.650 0.460 795.110 ;
    END
  END wd_in[336]
  PIN wd_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 795.110 0.460 795.570 ;
    END
  END wd_in[337]
  PIN wd_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 795.570 0.460 796.030 ;
    END
  END wd_in[338]
  PIN wd_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 796.030 0.460 796.490 ;
    END
  END wd_in[339]
  PIN wd_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 796.490 0.460 796.950 ;
    END
  END wd_in[340]
  PIN wd_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 796.950 0.460 797.410 ;
    END
  END wd_in[341]
  PIN wd_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 797.410 0.460 797.870 ;
    END
  END wd_in[342]
  PIN wd_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 797.870 0.460 798.330 ;
    END
  END wd_in[343]
  PIN wd_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 798.330 0.460 798.790 ;
    END
  END wd_in[344]
  PIN wd_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 798.790 0.460 799.250 ;
    END
  END wd_in[345]
  PIN wd_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 799.250 0.460 799.710 ;
    END
  END wd_in[346]
  PIN wd_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 799.710 0.460 800.170 ;
    END
  END wd_in[347]
  PIN wd_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 800.170 0.460 800.630 ;
    END
  END wd_in[348]
  PIN wd_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 800.630 0.460 801.090 ;
    END
  END wd_in[349]
  PIN wd_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 801.090 0.460 801.550 ;
    END
  END wd_in[350]
  PIN wd_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 801.550 0.460 802.010 ;
    END
  END wd_in[351]
  PIN wd_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 802.010 0.460 802.470 ;
    END
  END wd_in[352]
  PIN wd_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 802.470 0.460 802.930 ;
    END
  END wd_in[353]
  PIN wd_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 802.930 0.460 803.390 ;
    END
  END wd_in[354]
  PIN wd_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 803.390 0.460 803.850 ;
    END
  END wd_in[355]
  PIN wd_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 803.850 0.460 804.310 ;
    END
  END wd_in[356]
  PIN wd_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 804.310 0.460 804.770 ;
    END
  END wd_in[357]
  PIN wd_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 804.770 0.460 805.230 ;
    END
  END wd_in[358]
  PIN wd_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 805.230 0.460 805.690 ;
    END
  END wd_in[359]
  PIN wd_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 805.690 0.460 806.150 ;
    END
  END wd_in[360]
  PIN wd_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 806.150 0.460 806.610 ;
    END
  END wd_in[361]
  PIN wd_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 806.610 0.460 807.070 ;
    END
  END wd_in[362]
  PIN wd_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 807.070 0.460 807.530 ;
    END
  END wd_in[363]
  PIN wd_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 807.530 0.460 807.990 ;
    END
  END wd_in[364]
  PIN wd_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 807.990 0.460 808.450 ;
    END
  END wd_in[365]
  PIN wd_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 808.450 0.460 808.910 ;
    END
  END wd_in[366]
  PIN wd_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 808.910 0.460 809.370 ;
    END
  END wd_in[367]
  PIN wd_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 809.370 0.460 809.830 ;
    END
  END wd_in[368]
  PIN wd_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 809.830 0.460 810.290 ;
    END
  END wd_in[369]
  PIN wd_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 810.290 0.460 810.750 ;
    END
  END wd_in[370]
  PIN wd_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 810.750 0.460 811.210 ;
    END
  END wd_in[371]
  PIN wd_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 811.210 0.460 811.670 ;
    END
  END wd_in[372]
  PIN wd_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 811.670 0.460 812.130 ;
    END
  END wd_in[373]
  PIN wd_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 812.130 0.460 812.590 ;
    END
  END wd_in[374]
  PIN wd_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 812.590 0.460 813.050 ;
    END
  END wd_in[375]
  PIN wd_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 813.050 0.460 813.510 ;
    END
  END wd_in[376]
  PIN wd_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 813.510 0.460 813.970 ;
    END
  END wd_in[377]
  PIN wd_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 813.970 0.460 814.430 ;
    END
  END wd_in[378]
  PIN wd_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 814.430 0.460 814.890 ;
    END
  END wd_in[379]
  PIN wd_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 814.890 0.460 815.350 ;
    END
  END wd_in[380]
  PIN wd_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 815.350 0.460 815.810 ;
    END
  END wd_in[381]
  PIN wd_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 815.810 0.460 816.270 ;
    END
  END wd_in[382]
  PIN wd_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 816.270 0.460 816.730 ;
    END
  END wd_in[383]
  PIN wd_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 816.730 0.460 817.190 ;
    END
  END wd_in[384]
  PIN wd_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 817.190 0.460 817.650 ;
    END
  END wd_in[385]
  PIN wd_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 817.650 0.460 818.110 ;
    END
  END wd_in[386]
  PIN wd_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 818.110 0.460 818.570 ;
    END
  END wd_in[387]
  PIN wd_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 818.570 0.460 819.030 ;
    END
  END wd_in[388]
  PIN wd_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 819.030 0.460 819.490 ;
    END
  END wd_in[389]
  PIN wd_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 819.490 0.460 819.950 ;
    END
  END wd_in[390]
  PIN wd_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 819.950 0.460 820.410 ;
    END
  END wd_in[391]
  PIN wd_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 820.410 0.460 820.870 ;
    END
  END wd_in[392]
  PIN wd_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 820.870 0.460 821.330 ;
    END
  END wd_in[393]
  PIN wd_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 821.330 0.460 821.790 ;
    END
  END wd_in[394]
  PIN wd_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 821.790 0.460 822.250 ;
    END
  END wd_in[395]
  PIN wd_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 822.250 0.460 822.710 ;
    END
  END wd_in[396]
  PIN wd_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 822.710 0.460 823.170 ;
    END
  END wd_in[397]
  PIN wd_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 823.170 0.460 823.630 ;
    END
  END wd_in[398]
  PIN wd_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 823.630 0.460 824.090 ;
    END
  END wd_in[399]
  PIN wd_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 824.090 0.460 824.550 ;
    END
  END wd_in[400]
  PIN wd_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 824.550 0.460 825.010 ;
    END
  END wd_in[401]
  PIN wd_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 825.010 0.460 825.470 ;
    END
  END wd_in[402]
  PIN wd_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 825.470 0.460 825.930 ;
    END
  END wd_in[403]
  PIN wd_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 825.930 0.460 826.390 ;
    END
  END wd_in[404]
  PIN wd_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 826.390 0.460 826.850 ;
    END
  END wd_in[405]
  PIN wd_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 826.850 0.460 827.310 ;
    END
  END wd_in[406]
  PIN wd_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 827.310 0.460 827.770 ;
    END
  END wd_in[407]
  PIN wd_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 827.770 0.460 828.230 ;
    END
  END wd_in[408]
  PIN wd_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 828.230 0.460 828.690 ;
    END
  END wd_in[409]
  PIN wd_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 828.690 0.460 829.150 ;
    END
  END wd_in[410]
  PIN wd_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 829.150 0.460 829.610 ;
    END
  END wd_in[411]
  PIN wd_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 829.610 0.460 830.070 ;
    END
  END wd_in[412]
  PIN wd_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 830.070 0.460 830.530 ;
    END
  END wd_in[413]
  PIN wd_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 830.530 0.460 830.990 ;
    END
  END wd_in[414]
  PIN wd_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 830.990 0.460 831.450 ;
    END
  END wd_in[415]
  PIN wd_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 831.450 0.460 831.910 ;
    END
  END wd_in[416]
  PIN wd_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 831.910 0.460 832.370 ;
    END
  END wd_in[417]
  PIN wd_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 832.370 0.460 832.830 ;
    END
  END wd_in[418]
  PIN wd_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 832.830 0.460 833.290 ;
    END
  END wd_in[419]
  PIN wd_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 833.290 0.460 833.750 ;
    END
  END wd_in[420]
  PIN wd_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 833.750 0.460 834.210 ;
    END
  END wd_in[421]
  PIN wd_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 834.210 0.460 834.670 ;
    END
  END wd_in[422]
  PIN wd_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 834.670 0.460 835.130 ;
    END
  END wd_in[423]
  PIN wd_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 835.130 0.460 835.590 ;
    END
  END wd_in[424]
  PIN wd_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 835.590 0.460 836.050 ;
    END
  END wd_in[425]
  PIN wd_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 836.050 0.460 836.510 ;
    END
  END wd_in[426]
  PIN wd_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 836.510 0.460 836.970 ;
    END
  END wd_in[427]
  PIN wd_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 836.970 0.460 837.430 ;
    END
  END wd_in[428]
  PIN wd_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 837.430 0.460 837.890 ;
    END
  END wd_in[429]
  PIN wd_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 837.890 0.460 838.350 ;
    END
  END wd_in[430]
  PIN wd_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 838.350 0.460 838.810 ;
    END
  END wd_in[431]
  PIN wd_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 838.810 0.460 839.270 ;
    END
  END wd_in[432]
  PIN wd_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 839.270 0.460 839.730 ;
    END
  END wd_in[433]
  PIN wd_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 839.730 0.460 840.190 ;
    END
  END wd_in[434]
  PIN wd_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 840.190 0.460 840.650 ;
    END
  END wd_in[435]
  PIN wd_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 840.650 0.460 841.110 ;
    END
  END wd_in[436]
  PIN wd_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 841.110 0.460 841.570 ;
    END
  END wd_in[437]
  PIN wd_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 841.570 0.460 842.030 ;
    END
  END wd_in[438]
  PIN wd_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 842.030 0.460 842.490 ;
    END
  END wd_in[439]
  PIN wd_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 842.490 0.460 842.950 ;
    END
  END wd_in[440]
  PIN wd_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 842.950 0.460 843.410 ;
    END
  END wd_in[441]
  PIN wd_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 843.410 0.460 843.870 ;
    END
  END wd_in[442]
  PIN wd_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 843.870 0.460 844.330 ;
    END
  END wd_in[443]
  PIN wd_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 844.330 0.460 844.790 ;
    END
  END wd_in[444]
  PIN wd_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 844.790 0.460 845.250 ;
    END
  END wd_in[445]
  PIN wd_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 845.250 0.460 845.710 ;
    END
  END wd_in[446]
  PIN wd_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 845.710 0.460 846.170 ;
    END
  END wd_in[447]
  PIN wd_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 846.170 0.460 846.630 ;
    END
  END wd_in[448]
  PIN wd_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 846.630 0.460 847.090 ;
    END
  END wd_in[449]
  PIN wd_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 847.090 0.460 847.550 ;
    END
  END wd_in[450]
  PIN wd_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 847.550 0.460 848.010 ;
    END
  END wd_in[451]
  PIN wd_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 848.010 0.460 848.470 ;
    END
  END wd_in[452]
  PIN wd_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 848.470 0.460 848.930 ;
    END
  END wd_in[453]
  PIN wd_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 848.930 0.460 849.390 ;
    END
  END wd_in[454]
  PIN wd_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 849.390 0.460 849.850 ;
    END
  END wd_in[455]
  PIN wd_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 849.850 0.460 850.310 ;
    END
  END wd_in[456]
  PIN wd_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 850.310 0.460 850.770 ;
    END
  END wd_in[457]
  PIN wd_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 850.770 0.460 851.230 ;
    END
  END wd_in[458]
  PIN wd_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 851.230 0.460 851.690 ;
    END
  END wd_in[459]
  PIN wd_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 851.690 0.460 852.150 ;
    END
  END wd_in[460]
  PIN wd_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 852.150 0.460 852.610 ;
    END
  END wd_in[461]
  PIN wd_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 852.610 0.460 853.070 ;
    END
  END wd_in[462]
  PIN wd_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 853.070 0.460 853.530 ;
    END
  END wd_in[463]
  PIN wd_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 853.530 0.460 853.990 ;
    END
  END wd_in[464]
  PIN wd_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 853.990 0.460 854.450 ;
    END
  END wd_in[465]
  PIN wd_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 854.450 0.460 854.910 ;
    END
  END wd_in[466]
  PIN wd_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 854.910 0.460 855.370 ;
    END
  END wd_in[467]
  PIN wd_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 855.370 0.460 855.830 ;
    END
  END wd_in[468]
  PIN wd_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 855.830 0.460 856.290 ;
    END
  END wd_in[469]
  PIN wd_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 856.290 0.460 856.750 ;
    END
  END wd_in[470]
  PIN wd_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 856.750 0.460 857.210 ;
    END
  END wd_in[471]
  PIN wd_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 857.210 0.460 857.670 ;
    END
  END wd_in[472]
  PIN wd_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 857.670 0.460 858.130 ;
    END
  END wd_in[473]
  PIN wd_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 858.130 0.460 858.590 ;
    END
  END wd_in[474]
  PIN wd_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 858.590 0.460 859.050 ;
    END
  END wd_in[475]
  PIN wd_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 859.050 0.460 859.510 ;
    END
  END wd_in[476]
  PIN wd_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 859.510 0.460 859.970 ;
    END
  END wd_in[477]
  PIN wd_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 859.970 0.460 860.430 ;
    END
  END wd_in[478]
  PIN wd_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 860.430 0.460 860.890 ;
    END
  END wd_in[479]
  PIN wd_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 860.890 0.460 861.350 ;
    END
  END wd_in[480]
  PIN wd_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 861.350 0.460 861.810 ;
    END
  END wd_in[481]
  PIN wd_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 861.810 0.460 862.270 ;
    END
  END wd_in[482]
  PIN wd_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 862.270 0.460 862.730 ;
    END
  END wd_in[483]
  PIN wd_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 862.730 0.460 863.190 ;
    END
  END wd_in[484]
  PIN wd_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 863.190 0.460 863.650 ;
    END
  END wd_in[485]
  PIN wd_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 863.650 0.460 864.110 ;
    END
  END wd_in[486]
  PIN wd_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 864.110 0.460 864.570 ;
    END
  END wd_in[487]
  PIN wd_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 864.570 0.460 865.030 ;
    END
  END wd_in[488]
  PIN wd_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 865.030 0.460 865.490 ;
    END
  END wd_in[489]
  PIN wd_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 865.490 0.460 865.950 ;
    END
  END wd_in[490]
  PIN wd_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 865.950 0.460 866.410 ;
    END
  END wd_in[491]
  PIN wd_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 866.410 0.460 866.870 ;
    END
  END wd_in[492]
  PIN wd_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 866.870 0.460 867.330 ;
    END
  END wd_in[493]
  PIN wd_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 867.330 0.460 867.790 ;
    END
  END wd_in[494]
  PIN wd_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 867.790 0.460 868.250 ;
    END
  END wd_in[495]
  PIN wd_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 868.250 0.460 868.710 ;
    END
  END wd_in[496]
  PIN wd_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 868.710 0.460 869.170 ;
    END
  END wd_in[497]
  PIN wd_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 869.170 0.460 869.630 ;
    END
  END wd_in[498]
  PIN wd_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 869.630 0.460 870.090 ;
    END
  END wd_in[499]
  PIN wd_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 870.090 0.460 870.550 ;
    END
  END wd_in[500]
  PIN wd_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 870.550 0.460 871.010 ;
    END
  END wd_in[501]
  PIN wd_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 871.010 0.460 871.470 ;
    END
  END wd_in[502]
  PIN wd_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 871.470 0.460 871.930 ;
    END
  END wd_in[503]
  PIN wd_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 871.930 0.460 872.390 ;
    END
  END wd_in[504]
  PIN wd_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 872.390 0.460 872.850 ;
    END
  END wd_in[505]
  PIN wd_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 872.850 0.460 873.310 ;
    END
  END wd_in[506]
  PIN wd_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 873.310 0.460 873.770 ;
    END
  END wd_in[507]
  PIN wd_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 873.770 0.460 874.230 ;
    END
  END wd_in[508]
  PIN wd_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 874.230 0.460 874.690 ;
    END
  END wd_in[509]
  PIN wd_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 874.690 0.460 875.150 ;
    END
  END wd_in[510]
  PIN wd_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 875.150 0.460 875.610 ;
    END
  END wd_in[511]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 957.950 0.460 958.410 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 958.410 0.460 958.870 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 958.870 0.460 959.330 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 959.330 0.460 959.790 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 959.790 0.460 960.250 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 960.250 0.460 960.710 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 960.710 0.460 961.170 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 961.170 0.460 961.630 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1043.970 0.460 1044.430 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1044.430 0.460 1044.890 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1044.890 0.460 1045.350 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.680 4.600 5.520 1048.040 ;
      RECT 11.040 4.600 12.880 1048.040 ;
      RECT 18.400 4.600 20.240 1048.040 ;
      RECT 25.760 4.600 27.600 1048.040 ;
      RECT 33.120 4.600 34.960 1048.040 ;
      RECT 40.480 4.600 42.320 1048.040 ;
      RECT 47.840 4.600 49.680 1048.040 ;
      RECT 55.200 4.600 57.040 1048.040 ;
      RECT 62.560 4.600 64.400 1048.040 ;
      RECT 69.920 4.600 71.760 1048.040 ;
      RECT 77.280 4.600 79.120 1048.040 ;
      RECT 84.640 4.600 86.480 1048.040 ;
      RECT 92.000 4.600 93.840 1048.040 ;
      RECT 99.360 4.600 101.200 1048.040 ;
      RECT 106.720 4.600 108.560 1048.040 ;
      RECT 114.080 4.600 115.920 1048.040 ;
      RECT 121.440 4.600 123.280 1048.040 ;
      RECT 128.800 4.600 130.640 1048.040 ;
      RECT 136.160 4.600 138.000 1048.040 ;
      RECT 143.520 4.600 145.360 1048.040 ;
      RECT 150.880 4.600 152.720 1048.040 ;
      RECT 158.240 4.600 160.080 1048.040 ;
      RECT 165.600 4.600 167.440 1048.040 ;
      RECT 172.960 4.600 174.800 1048.040 ;
      RECT 180.320 4.600 182.160 1048.040 ;
      RECT 187.680 4.600 189.520 1048.040 ;
      RECT 195.040 4.600 196.880 1048.040 ;
      RECT 202.400 4.600 204.240 1048.040 ;
      RECT 209.760 4.600 211.600 1048.040 ;
      RECT 217.120 4.600 218.960 1048.040 ;
      RECT 224.480 4.600 226.320 1048.040 ;
      RECT 231.840 4.600 233.680 1048.040 ;
      RECT 239.200 4.600 241.040 1048.040 ;
      RECT 246.560 4.600 248.400 1048.040 ;
      RECT 253.920 4.600 255.760 1048.040 ;
      RECT 261.280 4.600 263.120 1048.040 ;
      RECT 268.640 4.600 270.480 1048.040 ;
      RECT 276.000 4.600 277.840 1048.040 ;
      RECT 283.360 4.600 285.200 1048.040 ;
      RECT 290.720 4.600 292.560 1048.040 ;
      RECT 298.080 4.600 299.920 1048.040 ;
      RECT 305.440 4.600 307.280 1048.040 ;
      RECT 312.800 4.600 314.640 1048.040 ;
      RECT 320.160 4.600 322.000 1048.040 ;
      RECT 327.520 4.600 329.360 1048.040 ;
      RECT 334.880 4.600 336.720 1048.040 ;
      RECT 342.240 4.600 344.080 1048.040 ;
      RECT 349.600 4.600 351.440 1048.040 ;
      RECT 356.960 4.600 358.800 1048.040 ;
      RECT 364.320 4.600 366.160 1048.040 ;
      RECT 371.680 4.600 373.520 1048.040 ;
      RECT 379.040 4.600 380.880 1048.040 ;
      RECT 386.400 4.600 388.240 1048.040 ;
      RECT 393.760 4.600 395.600 1048.040 ;
      RECT 401.120 4.600 402.960 1048.040 ;
      RECT 408.480 4.600 410.320 1048.040 ;
      RECT 415.840 4.600 417.680 1048.040 ;
      RECT 423.200 4.600 425.040 1048.040 ;
      RECT 430.560 4.600 432.400 1048.040 ;
      RECT 437.920 4.600 439.760 1048.040 ;
      RECT 445.280 4.600 447.120 1048.040 ;
      RECT 452.640 4.600 454.480 1048.040 ;
      RECT 460.000 4.600 461.840 1048.040 ;
      RECT 467.360 4.600 469.200 1048.040 ;
      RECT 474.720 4.600 476.560 1048.040 ;
      RECT 482.080 4.600 483.920 1048.040 ;
      RECT 489.440 4.600 491.280 1048.040 ;
      RECT 496.800 4.600 498.640 1048.040 ;
      RECT 504.160 4.600 506.000 1048.040 ;
      RECT 511.520 4.600 513.360 1048.040 ;
      RECT 518.880 4.600 520.720 1048.040 ;
      RECT 526.240 4.600 528.080 1048.040 ;
      RECT 533.600 4.600 535.440 1048.040 ;
      RECT 540.960 4.600 542.800 1048.040 ;
      RECT 548.320 4.600 550.160 1048.040 ;
      RECT 555.680 4.600 557.520 1048.040 ;
      RECT 563.040 4.600 564.880 1048.040 ;
      RECT 570.400 4.600 572.240 1048.040 ;
      RECT 577.760 4.600 579.600 1048.040 ;
      RECT 585.120 4.600 586.960 1048.040 ;
      RECT 592.480 4.600 594.320 1048.040 ;
      RECT 599.840 4.600 601.680 1048.040 ;
      RECT 607.200 4.600 609.040 1048.040 ;
      RECT 614.560 4.600 616.400 1048.040 ;
      RECT 621.920 4.600 623.760 1048.040 ;
      RECT 629.280 4.600 631.120 1048.040 ;
      RECT 636.640 4.600 638.480 1048.040 ;
      RECT 644.000 4.600 645.840 1048.040 ;
      RECT 651.360 4.600 653.200 1048.040 ;
      RECT 658.720 4.600 660.560 1048.040 ;
      RECT 666.080 4.600 667.920 1048.040 ;
      RECT 673.440 4.600 675.280 1048.040 ;
      RECT 680.800 4.600 682.640 1048.040 ;
      RECT 688.160 4.600 690.000 1048.040 ;
      RECT 695.520 4.600 697.360 1048.040 ;
      RECT 702.880 4.600 704.720 1048.040 ;
      RECT 710.240 4.600 712.080 1048.040 ;
      RECT 717.600 4.600 719.440 1048.040 ;
      RECT 724.960 4.600 726.800 1048.040 ;
      RECT 732.320 4.600 734.160 1048.040 ;
      RECT 739.680 4.600 741.520 1048.040 ;
      RECT 747.040 4.600 748.880 1048.040 ;
      RECT 754.400 4.600 756.240 1048.040 ;
      RECT 761.760 4.600 763.600 1048.040 ;
      RECT 769.120 4.600 770.960 1048.040 ;
      RECT 776.480 4.600 778.320 1048.040 ;
      RECT 783.840 4.600 785.680 1048.040 ;
      RECT 791.200 4.600 793.040 1048.040 ;
      RECT 798.560 4.600 800.400 1048.040 ;
      RECT 805.920 4.600 807.760 1048.040 ;
      RECT 813.280 4.600 815.120 1048.040 ;
      RECT 820.640 4.600 822.480 1048.040 ;
      RECT 828.000 4.600 829.840 1048.040 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 7.360 4.600 9.200 1048.040 ;
      RECT 14.720 4.600 16.560 1048.040 ;
      RECT 22.080 4.600 23.920 1048.040 ;
      RECT 29.440 4.600 31.280 1048.040 ;
      RECT 36.800 4.600 38.640 1048.040 ;
      RECT 44.160 4.600 46.000 1048.040 ;
      RECT 51.520 4.600 53.360 1048.040 ;
      RECT 58.880 4.600 60.720 1048.040 ;
      RECT 66.240 4.600 68.080 1048.040 ;
      RECT 73.600 4.600 75.440 1048.040 ;
      RECT 80.960 4.600 82.800 1048.040 ;
      RECT 88.320 4.600 90.160 1048.040 ;
      RECT 95.680 4.600 97.520 1048.040 ;
      RECT 103.040 4.600 104.880 1048.040 ;
      RECT 110.400 4.600 112.240 1048.040 ;
      RECT 117.760 4.600 119.600 1048.040 ;
      RECT 125.120 4.600 126.960 1048.040 ;
      RECT 132.480 4.600 134.320 1048.040 ;
      RECT 139.840 4.600 141.680 1048.040 ;
      RECT 147.200 4.600 149.040 1048.040 ;
      RECT 154.560 4.600 156.400 1048.040 ;
      RECT 161.920 4.600 163.760 1048.040 ;
      RECT 169.280 4.600 171.120 1048.040 ;
      RECT 176.640 4.600 178.480 1048.040 ;
      RECT 184.000 4.600 185.840 1048.040 ;
      RECT 191.360 4.600 193.200 1048.040 ;
      RECT 198.720 4.600 200.560 1048.040 ;
      RECT 206.080 4.600 207.920 1048.040 ;
      RECT 213.440 4.600 215.280 1048.040 ;
      RECT 220.800 4.600 222.640 1048.040 ;
      RECT 228.160 4.600 230.000 1048.040 ;
      RECT 235.520 4.600 237.360 1048.040 ;
      RECT 242.880 4.600 244.720 1048.040 ;
      RECT 250.240 4.600 252.080 1048.040 ;
      RECT 257.600 4.600 259.440 1048.040 ;
      RECT 264.960 4.600 266.800 1048.040 ;
      RECT 272.320 4.600 274.160 1048.040 ;
      RECT 279.680 4.600 281.520 1048.040 ;
      RECT 287.040 4.600 288.880 1048.040 ;
      RECT 294.400 4.600 296.240 1048.040 ;
      RECT 301.760 4.600 303.600 1048.040 ;
      RECT 309.120 4.600 310.960 1048.040 ;
      RECT 316.480 4.600 318.320 1048.040 ;
      RECT 323.840 4.600 325.680 1048.040 ;
      RECT 331.200 4.600 333.040 1048.040 ;
      RECT 338.560 4.600 340.400 1048.040 ;
      RECT 345.920 4.600 347.760 1048.040 ;
      RECT 353.280 4.600 355.120 1048.040 ;
      RECT 360.640 4.600 362.480 1048.040 ;
      RECT 368.000 4.600 369.840 1048.040 ;
      RECT 375.360 4.600 377.200 1048.040 ;
      RECT 382.720 4.600 384.560 1048.040 ;
      RECT 390.080 4.600 391.920 1048.040 ;
      RECT 397.440 4.600 399.280 1048.040 ;
      RECT 404.800 4.600 406.640 1048.040 ;
      RECT 412.160 4.600 414.000 1048.040 ;
      RECT 419.520 4.600 421.360 1048.040 ;
      RECT 426.880 4.600 428.720 1048.040 ;
      RECT 434.240 4.600 436.080 1048.040 ;
      RECT 441.600 4.600 443.440 1048.040 ;
      RECT 448.960 4.600 450.800 1048.040 ;
      RECT 456.320 4.600 458.160 1048.040 ;
      RECT 463.680 4.600 465.520 1048.040 ;
      RECT 471.040 4.600 472.880 1048.040 ;
      RECT 478.400 4.600 480.240 1048.040 ;
      RECT 485.760 4.600 487.600 1048.040 ;
      RECT 493.120 4.600 494.960 1048.040 ;
      RECT 500.480 4.600 502.320 1048.040 ;
      RECT 507.840 4.600 509.680 1048.040 ;
      RECT 515.200 4.600 517.040 1048.040 ;
      RECT 522.560 4.600 524.400 1048.040 ;
      RECT 529.920 4.600 531.760 1048.040 ;
      RECT 537.280 4.600 539.120 1048.040 ;
      RECT 544.640 4.600 546.480 1048.040 ;
      RECT 552.000 4.600 553.840 1048.040 ;
      RECT 559.360 4.600 561.200 1048.040 ;
      RECT 566.720 4.600 568.560 1048.040 ;
      RECT 574.080 4.600 575.920 1048.040 ;
      RECT 581.440 4.600 583.280 1048.040 ;
      RECT 588.800 4.600 590.640 1048.040 ;
      RECT 596.160 4.600 598.000 1048.040 ;
      RECT 603.520 4.600 605.360 1048.040 ;
      RECT 610.880 4.600 612.720 1048.040 ;
      RECT 618.240 4.600 620.080 1048.040 ;
      RECT 625.600 4.600 627.440 1048.040 ;
      RECT 632.960 4.600 634.800 1048.040 ;
      RECT 640.320 4.600 642.160 1048.040 ;
      RECT 647.680 4.600 649.520 1048.040 ;
      RECT 655.040 4.600 656.880 1048.040 ;
      RECT 662.400 4.600 664.240 1048.040 ;
      RECT 669.760 4.600 671.600 1048.040 ;
      RECT 677.120 4.600 678.960 1048.040 ;
      RECT 684.480 4.600 686.320 1048.040 ;
      RECT 691.840 4.600 693.680 1048.040 ;
      RECT 699.200 4.600 701.040 1048.040 ;
      RECT 706.560 4.600 708.400 1048.040 ;
      RECT 713.920 4.600 715.760 1048.040 ;
      RECT 721.280 4.600 723.120 1048.040 ;
      RECT 728.640 4.600 730.480 1048.040 ;
      RECT 736.000 4.600 737.840 1048.040 ;
      RECT 743.360 4.600 745.200 1048.040 ;
      RECT 750.720 4.600 752.560 1048.040 ;
      RECT 758.080 4.600 759.920 1048.040 ;
      RECT 765.440 4.600 767.280 1048.040 ;
      RECT 772.800 4.600 774.640 1048.040 ;
      RECT 780.160 4.600 782.000 1048.040 ;
      RECT 787.520 4.600 789.360 1048.040 ;
      RECT 794.880 4.600 796.720 1048.040 ;
      RECT 802.240 4.600 804.080 1048.040 ;
      RECT 809.600 4.600 811.440 1048.040 ;
      RECT 816.960 4.600 818.800 1048.040 ;
      RECT 824.320 4.600 826.160 1048.040 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 834.440 1052.640 ;
    LAYER met2 ;
    RECT 0 0 834.440 1052.640 ;
    LAYER met3 ;
    RECT 0.460 0 834.440 1052.640 ;
    RECT 0 0.000 0.460 4.370 ;
    RECT 0 4.830 0.460 4.830 ;
    RECT 0 5.290 0.460 5.290 ;
    RECT 0 5.750 0.460 5.750 ;
    RECT 0 6.210 0.460 6.210 ;
    RECT 0 6.670 0.460 6.670 ;
    RECT 0 7.130 0.460 7.130 ;
    RECT 0 7.590 0.460 7.590 ;
    RECT 0 8.050 0.460 8.050 ;
    RECT 0 8.510 0.460 8.510 ;
    RECT 0 8.970 0.460 8.970 ;
    RECT 0 9.430 0.460 9.430 ;
    RECT 0 9.890 0.460 9.890 ;
    RECT 0 10.350 0.460 10.350 ;
    RECT 0 10.810 0.460 10.810 ;
    RECT 0 11.270 0.460 11.270 ;
    RECT 0 11.730 0.460 11.730 ;
    RECT 0 12.190 0.460 12.190 ;
    RECT 0 12.650 0.460 12.650 ;
    RECT 0 13.110 0.460 13.110 ;
    RECT 0 13.570 0.460 13.570 ;
    RECT 0 14.030 0.460 14.030 ;
    RECT 0 14.490 0.460 14.490 ;
    RECT 0 14.950 0.460 14.950 ;
    RECT 0 15.410 0.460 15.410 ;
    RECT 0 15.870 0.460 15.870 ;
    RECT 0 16.330 0.460 16.330 ;
    RECT 0 16.790 0.460 16.790 ;
    RECT 0 17.250 0.460 17.250 ;
    RECT 0 17.710 0.460 17.710 ;
    RECT 0 18.170 0.460 18.170 ;
    RECT 0 18.630 0.460 18.630 ;
    RECT 0 19.090 0.460 19.090 ;
    RECT 0 19.550 0.460 19.550 ;
    RECT 0 20.010 0.460 20.010 ;
    RECT 0 20.470 0.460 20.470 ;
    RECT 0 20.930 0.460 20.930 ;
    RECT 0 21.390 0.460 21.390 ;
    RECT 0 21.850 0.460 21.850 ;
    RECT 0 22.310 0.460 22.310 ;
    RECT 0 22.770 0.460 22.770 ;
    RECT 0 23.230 0.460 23.230 ;
    RECT 0 23.690 0.460 23.690 ;
    RECT 0 24.150 0.460 24.150 ;
    RECT 0 24.610 0.460 24.610 ;
    RECT 0 25.070 0.460 25.070 ;
    RECT 0 25.530 0.460 25.530 ;
    RECT 0 25.990 0.460 25.990 ;
    RECT 0 26.450 0.460 26.450 ;
    RECT 0 26.910 0.460 26.910 ;
    RECT 0 27.370 0.460 27.370 ;
    RECT 0 27.830 0.460 27.830 ;
    RECT 0 28.290 0.460 28.290 ;
    RECT 0 28.750 0.460 28.750 ;
    RECT 0 29.210 0.460 29.210 ;
    RECT 0 29.670 0.460 29.670 ;
    RECT 0 30.130 0.460 30.130 ;
    RECT 0 30.590 0.460 30.590 ;
    RECT 0 31.050 0.460 31.050 ;
    RECT 0 31.510 0.460 31.510 ;
    RECT 0 31.970 0.460 31.970 ;
    RECT 0 32.430 0.460 32.430 ;
    RECT 0 32.890 0.460 32.890 ;
    RECT 0 33.350 0.460 33.350 ;
    RECT 0 33.810 0.460 33.810 ;
    RECT 0 34.270 0.460 34.270 ;
    RECT 0 34.730 0.460 34.730 ;
    RECT 0 35.190 0.460 35.190 ;
    RECT 0 35.650 0.460 35.650 ;
    RECT 0 36.110 0.460 36.110 ;
    RECT 0 36.570 0.460 36.570 ;
    RECT 0 37.030 0.460 37.030 ;
    RECT 0 37.490 0.460 37.490 ;
    RECT 0 37.950 0.460 37.950 ;
    RECT 0 38.410 0.460 38.410 ;
    RECT 0 38.870 0.460 38.870 ;
    RECT 0 39.330 0.460 39.330 ;
    RECT 0 39.790 0.460 39.790 ;
    RECT 0 40.250 0.460 40.250 ;
    RECT 0 40.710 0.460 40.710 ;
    RECT 0 41.170 0.460 41.170 ;
    RECT 0 41.630 0.460 41.630 ;
    RECT 0 42.090 0.460 42.090 ;
    RECT 0 42.550 0.460 42.550 ;
    RECT 0 43.010 0.460 43.010 ;
    RECT 0 43.470 0.460 43.470 ;
    RECT 0 43.930 0.460 43.930 ;
    RECT 0 44.390 0.460 44.390 ;
    RECT 0 44.850 0.460 44.850 ;
    RECT 0 45.310 0.460 45.310 ;
    RECT 0 45.770 0.460 45.770 ;
    RECT 0 46.230 0.460 46.230 ;
    RECT 0 46.690 0.460 46.690 ;
    RECT 0 47.150 0.460 47.150 ;
    RECT 0 47.610 0.460 47.610 ;
    RECT 0 48.070 0.460 48.070 ;
    RECT 0 48.530 0.460 48.530 ;
    RECT 0 48.990 0.460 48.990 ;
    RECT 0 49.450 0.460 49.450 ;
    RECT 0 49.910 0.460 49.910 ;
    RECT 0 50.370 0.460 50.370 ;
    RECT 0 50.830 0.460 50.830 ;
    RECT 0 51.290 0.460 51.290 ;
    RECT 0 51.750 0.460 51.750 ;
    RECT 0 52.210 0.460 52.210 ;
    RECT 0 52.670 0.460 52.670 ;
    RECT 0 53.130 0.460 53.130 ;
    RECT 0 53.590 0.460 53.590 ;
    RECT 0 54.050 0.460 54.050 ;
    RECT 0 54.510 0.460 54.510 ;
    RECT 0 54.970 0.460 54.970 ;
    RECT 0 55.430 0.460 55.430 ;
    RECT 0 55.890 0.460 55.890 ;
    RECT 0 56.350 0.460 56.350 ;
    RECT 0 56.810 0.460 56.810 ;
    RECT 0 57.270 0.460 57.270 ;
    RECT 0 57.730 0.460 57.730 ;
    RECT 0 58.190 0.460 58.190 ;
    RECT 0 58.650 0.460 58.650 ;
    RECT 0 59.110 0.460 59.110 ;
    RECT 0 59.570 0.460 59.570 ;
    RECT 0 60.030 0.460 60.030 ;
    RECT 0 60.490 0.460 60.490 ;
    RECT 0 60.950 0.460 60.950 ;
    RECT 0 61.410 0.460 61.410 ;
    RECT 0 61.870 0.460 61.870 ;
    RECT 0 62.330 0.460 62.330 ;
    RECT 0 62.790 0.460 62.790 ;
    RECT 0 63.250 0.460 63.250 ;
    RECT 0 63.710 0.460 63.710 ;
    RECT 0 64.170 0.460 64.170 ;
    RECT 0 64.630 0.460 64.630 ;
    RECT 0 65.090 0.460 65.090 ;
    RECT 0 65.550 0.460 65.550 ;
    RECT 0 66.010 0.460 66.010 ;
    RECT 0 66.470 0.460 66.470 ;
    RECT 0 66.930 0.460 66.930 ;
    RECT 0 67.390 0.460 67.390 ;
    RECT 0 67.850 0.460 67.850 ;
    RECT 0 68.310 0.460 68.310 ;
    RECT 0 68.770 0.460 68.770 ;
    RECT 0 69.230 0.460 69.230 ;
    RECT 0 69.690 0.460 69.690 ;
    RECT 0 70.150 0.460 70.150 ;
    RECT 0 70.610 0.460 70.610 ;
    RECT 0 71.070 0.460 71.070 ;
    RECT 0 71.530 0.460 71.530 ;
    RECT 0 71.990 0.460 71.990 ;
    RECT 0 72.450 0.460 72.450 ;
    RECT 0 72.910 0.460 72.910 ;
    RECT 0 73.370 0.460 73.370 ;
    RECT 0 73.830 0.460 73.830 ;
    RECT 0 74.290 0.460 74.290 ;
    RECT 0 74.750 0.460 74.750 ;
    RECT 0 75.210 0.460 75.210 ;
    RECT 0 75.670 0.460 75.670 ;
    RECT 0 76.130 0.460 76.130 ;
    RECT 0 76.590 0.460 76.590 ;
    RECT 0 77.050 0.460 77.050 ;
    RECT 0 77.510 0.460 77.510 ;
    RECT 0 77.970 0.460 77.970 ;
    RECT 0 78.430 0.460 78.430 ;
    RECT 0 78.890 0.460 78.890 ;
    RECT 0 79.350 0.460 79.350 ;
    RECT 0 79.810 0.460 79.810 ;
    RECT 0 80.270 0.460 80.270 ;
    RECT 0 80.730 0.460 80.730 ;
    RECT 0 81.190 0.460 81.190 ;
    RECT 0 81.650 0.460 81.650 ;
    RECT 0 82.110 0.460 82.110 ;
    RECT 0 82.570 0.460 82.570 ;
    RECT 0 83.030 0.460 83.030 ;
    RECT 0 83.490 0.460 83.490 ;
    RECT 0 83.950 0.460 83.950 ;
    RECT 0 84.410 0.460 84.410 ;
    RECT 0 84.870 0.460 84.870 ;
    RECT 0 85.330 0.460 85.330 ;
    RECT 0 85.790 0.460 85.790 ;
    RECT 0 86.250 0.460 86.250 ;
    RECT 0 86.710 0.460 86.710 ;
    RECT 0 87.170 0.460 87.170 ;
    RECT 0 87.630 0.460 87.630 ;
    RECT 0 88.090 0.460 88.090 ;
    RECT 0 88.550 0.460 88.550 ;
    RECT 0 89.010 0.460 89.010 ;
    RECT 0 89.470 0.460 89.470 ;
    RECT 0 89.930 0.460 89.930 ;
    RECT 0 90.390 0.460 90.390 ;
    RECT 0 90.850 0.460 90.850 ;
    RECT 0 91.310 0.460 91.310 ;
    RECT 0 91.770 0.460 91.770 ;
    RECT 0 92.230 0.460 92.230 ;
    RECT 0 92.690 0.460 92.690 ;
    RECT 0 93.150 0.460 93.150 ;
    RECT 0 93.610 0.460 93.610 ;
    RECT 0 94.070 0.460 94.070 ;
    RECT 0 94.530 0.460 94.530 ;
    RECT 0 94.990 0.460 94.990 ;
    RECT 0 95.450 0.460 95.450 ;
    RECT 0 95.910 0.460 95.910 ;
    RECT 0 96.370 0.460 96.370 ;
    RECT 0 96.830 0.460 96.830 ;
    RECT 0 97.290 0.460 97.290 ;
    RECT 0 97.750 0.460 97.750 ;
    RECT 0 98.210 0.460 98.210 ;
    RECT 0 98.670 0.460 98.670 ;
    RECT 0 99.130 0.460 99.130 ;
    RECT 0 99.590 0.460 99.590 ;
    RECT 0 100.050 0.460 100.050 ;
    RECT 0 100.510 0.460 100.510 ;
    RECT 0 100.970 0.460 100.970 ;
    RECT 0 101.430 0.460 101.430 ;
    RECT 0 101.890 0.460 101.890 ;
    RECT 0 102.350 0.460 102.350 ;
    RECT 0 102.810 0.460 102.810 ;
    RECT 0 103.270 0.460 103.270 ;
    RECT 0 103.730 0.460 103.730 ;
    RECT 0 104.190 0.460 104.190 ;
    RECT 0 104.650 0.460 104.650 ;
    RECT 0 105.110 0.460 105.110 ;
    RECT 0 105.570 0.460 105.570 ;
    RECT 0 106.030 0.460 106.030 ;
    RECT 0 106.490 0.460 106.490 ;
    RECT 0 106.950 0.460 106.950 ;
    RECT 0 107.410 0.460 107.410 ;
    RECT 0 107.870 0.460 107.870 ;
    RECT 0 108.330 0.460 108.330 ;
    RECT 0 108.790 0.460 108.790 ;
    RECT 0 109.250 0.460 109.250 ;
    RECT 0 109.710 0.460 109.710 ;
    RECT 0 110.170 0.460 110.170 ;
    RECT 0 110.630 0.460 110.630 ;
    RECT 0 111.090 0.460 111.090 ;
    RECT 0 111.550 0.460 111.550 ;
    RECT 0 112.010 0.460 112.010 ;
    RECT 0 112.470 0.460 112.470 ;
    RECT 0 112.930 0.460 112.930 ;
    RECT 0 113.390 0.460 113.390 ;
    RECT 0 113.850 0.460 113.850 ;
    RECT 0 114.310 0.460 114.310 ;
    RECT 0 114.770 0.460 114.770 ;
    RECT 0 115.230 0.460 115.230 ;
    RECT 0 115.690 0.460 115.690 ;
    RECT 0 116.150 0.460 116.150 ;
    RECT 0 116.610 0.460 116.610 ;
    RECT 0 117.070 0.460 117.070 ;
    RECT 0 117.530 0.460 117.530 ;
    RECT 0 117.990 0.460 117.990 ;
    RECT 0 118.450 0.460 118.450 ;
    RECT 0 118.910 0.460 118.910 ;
    RECT 0 119.370 0.460 119.370 ;
    RECT 0 119.830 0.460 119.830 ;
    RECT 0 120.290 0.460 120.290 ;
    RECT 0 120.750 0.460 120.750 ;
    RECT 0 121.210 0.460 121.210 ;
    RECT 0 121.670 0.460 121.670 ;
    RECT 0 122.130 0.460 122.130 ;
    RECT 0 122.590 0.460 122.590 ;
    RECT 0 123.050 0.460 123.050 ;
    RECT 0 123.510 0.460 123.510 ;
    RECT 0 123.970 0.460 123.970 ;
    RECT 0 124.430 0.460 124.430 ;
    RECT 0 124.890 0.460 124.890 ;
    RECT 0 125.350 0.460 125.350 ;
    RECT 0 125.810 0.460 125.810 ;
    RECT 0 126.270 0.460 126.270 ;
    RECT 0 126.730 0.460 126.730 ;
    RECT 0 127.190 0.460 127.190 ;
    RECT 0 127.650 0.460 127.650 ;
    RECT 0 128.110 0.460 128.110 ;
    RECT 0 128.570 0.460 128.570 ;
    RECT 0 129.030 0.460 129.030 ;
    RECT 0 129.490 0.460 129.490 ;
    RECT 0 129.950 0.460 129.950 ;
    RECT 0 130.410 0.460 130.410 ;
    RECT 0 130.870 0.460 130.870 ;
    RECT 0 131.330 0.460 131.330 ;
    RECT 0 131.790 0.460 131.790 ;
    RECT 0 132.250 0.460 132.250 ;
    RECT 0 132.710 0.460 132.710 ;
    RECT 0 133.170 0.460 133.170 ;
    RECT 0 133.630 0.460 133.630 ;
    RECT 0 134.090 0.460 134.090 ;
    RECT 0 134.550 0.460 134.550 ;
    RECT 0 135.010 0.460 135.010 ;
    RECT 0 135.470 0.460 135.470 ;
    RECT 0 135.930 0.460 135.930 ;
    RECT 0 136.390 0.460 136.390 ;
    RECT 0 136.850 0.460 136.850 ;
    RECT 0 137.310 0.460 137.310 ;
    RECT 0 137.770 0.460 137.770 ;
    RECT 0 138.230 0.460 138.230 ;
    RECT 0 138.690 0.460 138.690 ;
    RECT 0 139.150 0.460 139.150 ;
    RECT 0 139.610 0.460 139.610 ;
    RECT 0 140.070 0.460 140.070 ;
    RECT 0 140.530 0.460 140.530 ;
    RECT 0 140.990 0.460 140.990 ;
    RECT 0 141.450 0.460 141.450 ;
    RECT 0 141.910 0.460 141.910 ;
    RECT 0 142.370 0.460 142.370 ;
    RECT 0 142.830 0.460 142.830 ;
    RECT 0 143.290 0.460 143.290 ;
    RECT 0 143.750 0.460 143.750 ;
    RECT 0 144.210 0.460 144.210 ;
    RECT 0 144.670 0.460 144.670 ;
    RECT 0 145.130 0.460 145.130 ;
    RECT 0 145.590 0.460 145.590 ;
    RECT 0 146.050 0.460 146.050 ;
    RECT 0 146.510 0.460 146.510 ;
    RECT 0 146.970 0.460 146.970 ;
    RECT 0 147.430 0.460 147.430 ;
    RECT 0 147.890 0.460 147.890 ;
    RECT 0 148.350 0.460 148.350 ;
    RECT 0 148.810 0.460 148.810 ;
    RECT 0 149.270 0.460 149.270 ;
    RECT 0 149.730 0.460 149.730 ;
    RECT 0 150.190 0.460 150.190 ;
    RECT 0 150.650 0.460 150.650 ;
    RECT 0 151.110 0.460 151.110 ;
    RECT 0 151.570 0.460 151.570 ;
    RECT 0 152.030 0.460 152.030 ;
    RECT 0 152.490 0.460 152.490 ;
    RECT 0 152.950 0.460 152.950 ;
    RECT 0 153.410 0.460 153.410 ;
    RECT 0 153.870 0.460 153.870 ;
    RECT 0 154.330 0.460 154.330 ;
    RECT 0 154.790 0.460 154.790 ;
    RECT 0 155.250 0.460 155.250 ;
    RECT 0 155.710 0.460 155.710 ;
    RECT 0 156.170 0.460 156.170 ;
    RECT 0 156.630 0.460 156.630 ;
    RECT 0 157.090 0.460 157.090 ;
    RECT 0 157.550 0.460 157.550 ;
    RECT 0 158.010 0.460 158.010 ;
    RECT 0 158.470 0.460 158.470 ;
    RECT 0 158.930 0.460 158.930 ;
    RECT 0 159.390 0.460 159.390 ;
    RECT 0 159.850 0.460 159.850 ;
    RECT 0 160.310 0.460 160.310 ;
    RECT 0 160.770 0.460 160.770 ;
    RECT 0 161.230 0.460 161.230 ;
    RECT 0 161.690 0.460 161.690 ;
    RECT 0 162.150 0.460 162.150 ;
    RECT 0 162.610 0.460 162.610 ;
    RECT 0 163.070 0.460 163.070 ;
    RECT 0 163.530 0.460 163.530 ;
    RECT 0 163.990 0.460 163.990 ;
    RECT 0 164.450 0.460 164.450 ;
    RECT 0 164.910 0.460 164.910 ;
    RECT 0 165.370 0.460 165.370 ;
    RECT 0 165.830 0.460 165.830 ;
    RECT 0 166.290 0.460 166.290 ;
    RECT 0 166.750 0.460 166.750 ;
    RECT 0 167.210 0.460 167.210 ;
    RECT 0 167.670 0.460 167.670 ;
    RECT 0 168.130 0.460 168.130 ;
    RECT 0 168.590 0.460 168.590 ;
    RECT 0 169.050 0.460 169.050 ;
    RECT 0 169.510 0.460 169.510 ;
    RECT 0 169.970 0.460 169.970 ;
    RECT 0 170.430 0.460 170.430 ;
    RECT 0 170.890 0.460 170.890 ;
    RECT 0 171.350 0.460 171.350 ;
    RECT 0 171.810 0.460 171.810 ;
    RECT 0 172.270 0.460 172.270 ;
    RECT 0 172.730 0.460 172.730 ;
    RECT 0 173.190 0.460 173.190 ;
    RECT 0 173.650 0.460 173.650 ;
    RECT 0 174.110 0.460 174.110 ;
    RECT 0 174.570 0.460 174.570 ;
    RECT 0 175.030 0.460 175.030 ;
    RECT 0 175.490 0.460 175.490 ;
    RECT 0 175.950 0.460 175.950 ;
    RECT 0 176.410 0.460 176.410 ;
    RECT 0 176.870 0.460 176.870 ;
    RECT 0 177.330 0.460 177.330 ;
    RECT 0 177.790 0.460 177.790 ;
    RECT 0 178.250 0.460 178.250 ;
    RECT 0 178.710 0.460 178.710 ;
    RECT 0 179.170 0.460 179.170 ;
    RECT 0 179.630 0.460 179.630 ;
    RECT 0 180.090 0.460 180.090 ;
    RECT 0 180.550 0.460 180.550 ;
    RECT 0 181.010 0.460 181.010 ;
    RECT 0 181.470 0.460 181.470 ;
    RECT 0 181.930 0.460 181.930 ;
    RECT 0 182.390 0.460 182.390 ;
    RECT 0 182.850 0.460 182.850 ;
    RECT 0 183.310 0.460 183.310 ;
    RECT 0 183.770 0.460 183.770 ;
    RECT 0 184.230 0.460 184.230 ;
    RECT 0 184.690 0.460 184.690 ;
    RECT 0 185.150 0.460 185.150 ;
    RECT 0 185.610 0.460 185.610 ;
    RECT 0 186.070 0.460 186.070 ;
    RECT 0 186.530 0.460 186.530 ;
    RECT 0 186.990 0.460 186.990 ;
    RECT 0 187.450 0.460 187.450 ;
    RECT 0 187.910 0.460 187.910 ;
    RECT 0 188.370 0.460 188.370 ;
    RECT 0 188.830 0.460 188.830 ;
    RECT 0 189.290 0.460 189.290 ;
    RECT 0 189.750 0.460 189.750 ;
    RECT 0 190.210 0.460 190.210 ;
    RECT 0 190.670 0.460 190.670 ;
    RECT 0 191.130 0.460 191.130 ;
    RECT 0 191.590 0.460 191.590 ;
    RECT 0 192.050 0.460 192.050 ;
    RECT 0 192.510 0.460 192.510 ;
    RECT 0 192.970 0.460 192.970 ;
    RECT 0 193.430 0.460 193.430 ;
    RECT 0 193.890 0.460 193.890 ;
    RECT 0 194.350 0.460 194.350 ;
    RECT 0 194.810 0.460 194.810 ;
    RECT 0 195.270 0.460 195.270 ;
    RECT 0 195.730 0.460 195.730 ;
    RECT 0 196.190 0.460 196.190 ;
    RECT 0 196.650 0.460 196.650 ;
    RECT 0 197.110 0.460 197.110 ;
    RECT 0 197.570 0.460 197.570 ;
    RECT 0 198.030 0.460 198.030 ;
    RECT 0 198.490 0.460 198.490 ;
    RECT 0 198.950 0.460 198.950 ;
    RECT 0 199.410 0.460 199.410 ;
    RECT 0 199.870 0.460 199.870 ;
    RECT 0 200.330 0.460 200.330 ;
    RECT 0 200.790 0.460 200.790 ;
    RECT 0 201.250 0.460 201.250 ;
    RECT 0 201.710 0.460 201.710 ;
    RECT 0 202.170 0.460 202.170 ;
    RECT 0 202.630 0.460 202.630 ;
    RECT 0 203.090 0.460 203.090 ;
    RECT 0 203.550 0.460 203.550 ;
    RECT 0 204.010 0.460 204.010 ;
    RECT 0 204.470 0.460 204.470 ;
    RECT 0 204.930 0.460 204.930 ;
    RECT 0 205.390 0.460 205.390 ;
    RECT 0 205.850 0.460 205.850 ;
    RECT 0 206.310 0.460 206.310 ;
    RECT 0 206.770 0.460 206.770 ;
    RECT 0 207.230 0.460 207.230 ;
    RECT 0 207.690 0.460 207.690 ;
    RECT 0 208.150 0.460 208.150 ;
    RECT 0 208.610 0.460 208.610 ;
    RECT 0 209.070 0.460 209.070 ;
    RECT 0 209.530 0.460 209.530 ;
    RECT 0 209.990 0.460 209.990 ;
    RECT 0 210.450 0.460 210.450 ;
    RECT 0 210.910 0.460 210.910 ;
    RECT 0 211.370 0.460 211.370 ;
    RECT 0 211.830 0.460 211.830 ;
    RECT 0 212.290 0.460 212.290 ;
    RECT 0 212.750 0.460 212.750 ;
    RECT 0 213.210 0.460 213.210 ;
    RECT 0 213.670 0.460 213.670 ;
    RECT 0 214.130 0.460 214.130 ;
    RECT 0 214.590 0.460 214.590 ;
    RECT 0 215.050 0.460 215.050 ;
    RECT 0 215.510 0.460 215.510 ;
    RECT 0 215.970 0.460 215.970 ;
    RECT 0 216.430 0.460 216.430 ;
    RECT 0 216.890 0.460 216.890 ;
    RECT 0 217.350 0.460 217.350 ;
    RECT 0 217.810 0.460 217.810 ;
    RECT 0 218.270 0.460 218.270 ;
    RECT 0 218.730 0.460 218.730 ;
    RECT 0 219.190 0.460 219.190 ;
    RECT 0 219.650 0.460 219.650 ;
    RECT 0 220.110 0.460 220.110 ;
    RECT 0 220.570 0.460 220.570 ;
    RECT 0 221.030 0.460 221.030 ;
    RECT 0 221.490 0.460 221.490 ;
    RECT 0 221.950 0.460 221.950 ;
    RECT 0 222.410 0.460 222.410 ;
    RECT 0 222.870 0.460 222.870 ;
    RECT 0 223.330 0.460 223.330 ;
    RECT 0 223.790 0.460 223.790 ;
    RECT 0 224.250 0.460 224.250 ;
    RECT 0 224.710 0.460 224.710 ;
    RECT 0 225.170 0.460 225.170 ;
    RECT 0 225.630 0.460 225.630 ;
    RECT 0 226.090 0.460 226.090 ;
    RECT 0 226.550 0.460 226.550 ;
    RECT 0 227.010 0.460 227.010 ;
    RECT 0 227.470 0.460 227.470 ;
    RECT 0 227.930 0.460 227.930 ;
    RECT 0 228.390 0.460 228.390 ;
    RECT 0 228.850 0.460 228.850 ;
    RECT 0 229.310 0.460 229.310 ;
    RECT 0 229.770 0.460 229.770 ;
    RECT 0 230.230 0.460 230.230 ;
    RECT 0 230.690 0.460 230.690 ;
    RECT 0 231.150 0.460 231.150 ;
    RECT 0 231.610 0.460 231.610 ;
    RECT 0 232.070 0.460 232.070 ;
    RECT 0 232.530 0.460 232.530 ;
    RECT 0 232.990 0.460 232.990 ;
    RECT 0 233.450 0.460 233.450 ;
    RECT 0 233.910 0.460 233.910 ;
    RECT 0 234.370 0.460 234.370 ;
    RECT 0 234.830 0.460 234.830 ;
    RECT 0 235.290 0.460 235.290 ;
    RECT 0 235.750 0.460 235.750 ;
    RECT 0 236.210 0.460 236.210 ;
    RECT 0 236.670 0.460 236.670 ;
    RECT 0 237.130 0.460 237.130 ;
    RECT 0 237.590 0.460 237.590 ;
    RECT 0 238.050 0.460 238.050 ;
    RECT 0 238.510 0.460 238.510 ;
    RECT 0 238.970 0.460 238.970 ;
    RECT 0 239.430 0.460 239.430 ;
    RECT 0 239.890 0.460 322.230 ;
    RECT 0 322.690 0.460 322.690 ;
    RECT 0 323.150 0.460 323.150 ;
    RECT 0 323.610 0.460 323.610 ;
    RECT 0 324.070 0.460 324.070 ;
    RECT 0 324.530 0.460 324.530 ;
    RECT 0 324.990 0.460 324.990 ;
    RECT 0 325.450 0.460 325.450 ;
    RECT 0 325.910 0.460 325.910 ;
    RECT 0 326.370 0.460 326.370 ;
    RECT 0 326.830 0.460 326.830 ;
    RECT 0 327.290 0.460 327.290 ;
    RECT 0 327.750 0.460 327.750 ;
    RECT 0 328.210 0.460 328.210 ;
    RECT 0 328.670 0.460 328.670 ;
    RECT 0 329.130 0.460 329.130 ;
    RECT 0 329.590 0.460 329.590 ;
    RECT 0 330.050 0.460 330.050 ;
    RECT 0 330.510 0.460 330.510 ;
    RECT 0 330.970 0.460 330.970 ;
    RECT 0 331.430 0.460 331.430 ;
    RECT 0 331.890 0.460 331.890 ;
    RECT 0 332.350 0.460 332.350 ;
    RECT 0 332.810 0.460 332.810 ;
    RECT 0 333.270 0.460 333.270 ;
    RECT 0 333.730 0.460 333.730 ;
    RECT 0 334.190 0.460 334.190 ;
    RECT 0 334.650 0.460 334.650 ;
    RECT 0 335.110 0.460 335.110 ;
    RECT 0 335.570 0.460 335.570 ;
    RECT 0 336.030 0.460 336.030 ;
    RECT 0 336.490 0.460 336.490 ;
    RECT 0 336.950 0.460 336.950 ;
    RECT 0 337.410 0.460 337.410 ;
    RECT 0 337.870 0.460 337.870 ;
    RECT 0 338.330 0.460 338.330 ;
    RECT 0 338.790 0.460 338.790 ;
    RECT 0 339.250 0.460 339.250 ;
    RECT 0 339.710 0.460 339.710 ;
    RECT 0 340.170 0.460 340.170 ;
    RECT 0 340.630 0.460 340.630 ;
    RECT 0 341.090 0.460 341.090 ;
    RECT 0 341.550 0.460 341.550 ;
    RECT 0 342.010 0.460 342.010 ;
    RECT 0 342.470 0.460 342.470 ;
    RECT 0 342.930 0.460 342.930 ;
    RECT 0 343.390 0.460 343.390 ;
    RECT 0 343.850 0.460 343.850 ;
    RECT 0 344.310 0.460 344.310 ;
    RECT 0 344.770 0.460 344.770 ;
    RECT 0 345.230 0.460 345.230 ;
    RECT 0 345.690 0.460 345.690 ;
    RECT 0 346.150 0.460 346.150 ;
    RECT 0 346.610 0.460 346.610 ;
    RECT 0 347.070 0.460 347.070 ;
    RECT 0 347.530 0.460 347.530 ;
    RECT 0 347.990 0.460 347.990 ;
    RECT 0 348.450 0.460 348.450 ;
    RECT 0 348.910 0.460 348.910 ;
    RECT 0 349.370 0.460 349.370 ;
    RECT 0 349.830 0.460 349.830 ;
    RECT 0 350.290 0.460 350.290 ;
    RECT 0 350.750 0.460 350.750 ;
    RECT 0 351.210 0.460 351.210 ;
    RECT 0 351.670 0.460 351.670 ;
    RECT 0 352.130 0.460 352.130 ;
    RECT 0 352.590 0.460 352.590 ;
    RECT 0 353.050 0.460 353.050 ;
    RECT 0 353.510 0.460 353.510 ;
    RECT 0 353.970 0.460 353.970 ;
    RECT 0 354.430 0.460 354.430 ;
    RECT 0 354.890 0.460 354.890 ;
    RECT 0 355.350 0.460 355.350 ;
    RECT 0 355.810 0.460 355.810 ;
    RECT 0 356.270 0.460 356.270 ;
    RECT 0 356.730 0.460 356.730 ;
    RECT 0 357.190 0.460 357.190 ;
    RECT 0 357.650 0.460 357.650 ;
    RECT 0 358.110 0.460 358.110 ;
    RECT 0 358.570 0.460 358.570 ;
    RECT 0 359.030 0.460 359.030 ;
    RECT 0 359.490 0.460 359.490 ;
    RECT 0 359.950 0.460 359.950 ;
    RECT 0 360.410 0.460 360.410 ;
    RECT 0 360.870 0.460 360.870 ;
    RECT 0 361.330 0.460 361.330 ;
    RECT 0 361.790 0.460 361.790 ;
    RECT 0 362.250 0.460 362.250 ;
    RECT 0 362.710 0.460 362.710 ;
    RECT 0 363.170 0.460 363.170 ;
    RECT 0 363.630 0.460 363.630 ;
    RECT 0 364.090 0.460 364.090 ;
    RECT 0 364.550 0.460 364.550 ;
    RECT 0 365.010 0.460 365.010 ;
    RECT 0 365.470 0.460 365.470 ;
    RECT 0 365.930 0.460 365.930 ;
    RECT 0 366.390 0.460 366.390 ;
    RECT 0 366.850 0.460 366.850 ;
    RECT 0 367.310 0.460 367.310 ;
    RECT 0 367.770 0.460 367.770 ;
    RECT 0 368.230 0.460 368.230 ;
    RECT 0 368.690 0.460 368.690 ;
    RECT 0 369.150 0.460 369.150 ;
    RECT 0 369.610 0.460 369.610 ;
    RECT 0 370.070 0.460 370.070 ;
    RECT 0 370.530 0.460 370.530 ;
    RECT 0 370.990 0.460 370.990 ;
    RECT 0 371.450 0.460 371.450 ;
    RECT 0 371.910 0.460 371.910 ;
    RECT 0 372.370 0.460 372.370 ;
    RECT 0 372.830 0.460 372.830 ;
    RECT 0 373.290 0.460 373.290 ;
    RECT 0 373.750 0.460 373.750 ;
    RECT 0 374.210 0.460 374.210 ;
    RECT 0 374.670 0.460 374.670 ;
    RECT 0 375.130 0.460 375.130 ;
    RECT 0 375.590 0.460 375.590 ;
    RECT 0 376.050 0.460 376.050 ;
    RECT 0 376.510 0.460 376.510 ;
    RECT 0 376.970 0.460 376.970 ;
    RECT 0 377.430 0.460 377.430 ;
    RECT 0 377.890 0.460 377.890 ;
    RECT 0 378.350 0.460 378.350 ;
    RECT 0 378.810 0.460 378.810 ;
    RECT 0 379.270 0.460 379.270 ;
    RECT 0 379.730 0.460 379.730 ;
    RECT 0 380.190 0.460 380.190 ;
    RECT 0 380.650 0.460 380.650 ;
    RECT 0 381.110 0.460 381.110 ;
    RECT 0 381.570 0.460 381.570 ;
    RECT 0 382.030 0.460 382.030 ;
    RECT 0 382.490 0.460 382.490 ;
    RECT 0 382.950 0.460 382.950 ;
    RECT 0 383.410 0.460 383.410 ;
    RECT 0 383.870 0.460 383.870 ;
    RECT 0 384.330 0.460 384.330 ;
    RECT 0 384.790 0.460 384.790 ;
    RECT 0 385.250 0.460 385.250 ;
    RECT 0 385.710 0.460 385.710 ;
    RECT 0 386.170 0.460 386.170 ;
    RECT 0 386.630 0.460 386.630 ;
    RECT 0 387.090 0.460 387.090 ;
    RECT 0 387.550 0.460 387.550 ;
    RECT 0 388.010 0.460 388.010 ;
    RECT 0 388.470 0.460 388.470 ;
    RECT 0 388.930 0.460 388.930 ;
    RECT 0 389.390 0.460 389.390 ;
    RECT 0 389.850 0.460 389.850 ;
    RECT 0 390.310 0.460 390.310 ;
    RECT 0 390.770 0.460 390.770 ;
    RECT 0 391.230 0.460 391.230 ;
    RECT 0 391.690 0.460 391.690 ;
    RECT 0 392.150 0.460 392.150 ;
    RECT 0 392.610 0.460 392.610 ;
    RECT 0 393.070 0.460 393.070 ;
    RECT 0 393.530 0.460 393.530 ;
    RECT 0 393.990 0.460 393.990 ;
    RECT 0 394.450 0.460 394.450 ;
    RECT 0 394.910 0.460 394.910 ;
    RECT 0 395.370 0.460 395.370 ;
    RECT 0 395.830 0.460 395.830 ;
    RECT 0 396.290 0.460 396.290 ;
    RECT 0 396.750 0.460 396.750 ;
    RECT 0 397.210 0.460 397.210 ;
    RECT 0 397.670 0.460 397.670 ;
    RECT 0 398.130 0.460 398.130 ;
    RECT 0 398.590 0.460 398.590 ;
    RECT 0 399.050 0.460 399.050 ;
    RECT 0 399.510 0.460 399.510 ;
    RECT 0 399.970 0.460 399.970 ;
    RECT 0 400.430 0.460 400.430 ;
    RECT 0 400.890 0.460 400.890 ;
    RECT 0 401.350 0.460 401.350 ;
    RECT 0 401.810 0.460 401.810 ;
    RECT 0 402.270 0.460 402.270 ;
    RECT 0 402.730 0.460 402.730 ;
    RECT 0 403.190 0.460 403.190 ;
    RECT 0 403.650 0.460 403.650 ;
    RECT 0 404.110 0.460 404.110 ;
    RECT 0 404.570 0.460 404.570 ;
    RECT 0 405.030 0.460 405.030 ;
    RECT 0 405.490 0.460 405.490 ;
    RECT 0 405.950 0.460 405.950 ;
    RECT 0 406.410 0.460 406.410 ;
    RECT 0 406.870 0.460 406.870 ;
    RECT 0 407.330 0.460 407.330 ;
    RECT 0 407.790 0.460 407.790 ;
    RECT 0 408.250 0.460 408.250 ;
    RECT 0 408.710 0.460 408.710 ;
    RECT 0 409.170 0.460 409.170 ;
    RECT 0 409.630 0.460 409.630 ;
    RECT 0 410.090 0.460 410.090 ;
    RECT 0 410.550 0.460 410.550 ;
    RECT 0 411.010 0.460 411.010 ;
    RECT 0 411.470 0.460 411.470 ;
    RECT 0 411.930 0.460 411.930 ;
    RECT 0 412.390 0.460 412.390 ;
    RECT 0 412.850 0.460 412.850 ;
    RECT 0 413.310 0.460 413.310 ;
    RECT 0 413.770 0.460 413.770 ;
    RECT 0 414.230 0.460 414.230 ;
    RECT 0 414.690 0.460 414.690 ;
    RECT 0 415.150 0.460 415.150 ;
    RECT 0 415.610 0.460 415.610 ;
    RECT 0 416.070 0.460 416.070 ;
    RECT 0 416.530 0.460 416.530 ;
    RECT 0 416.990 0.460 416.990 ;
    RECT 0 417.450 0.460 417.450 ;
    RECT 0 417.910 0.460 417.910 ;
    RECT 0 418.370 0.460 418.370 ;
    RECT 0 418.830 0.460 418.830 ;
    RECT 0 419.290 0.460 419.290 ;
    RECT 0 419.750 0.460 419.750 ;
    RECT 0 420.210 0.460 420.210 ;
    RECT 0 420.670 0.460 420.670 ;
    RECT 0 421.130 0.460 421.130 ;
    RECT 0 421.590 0.460 421.590 ;
    RECT 0 422.050 0.460 422.050 ;
    RECT 0 422.510 0.460 422.510 ;
    RECT 0 422.970 0.460 422.970 ;
    RECT 0 423.430 0.460 423.430 ;
    RECT 0 423.890 0.460 423.890 ;
    RECT 0 424.350 0.460 424.350 ;
    RECT 0 424.810 0.460 424.810 ;
    RECT 0 425.270 0.460 425.270 ;
    RECT 0 425.730 0.460 425.730 ;
    RECT 0 426.190 0.460 426.190 ;
    RECT 0 426.650 0.460 426.650 ;
    RECT 0 427.110 0.460 427.110 ;
    RECT 0 427.570 0.460 427.570 ;
    RECT 0 428.030 0.460 428.030 ;
    RECT 0 428.490 0.460 428.490 ;
    RECT 0 428.950 0.460 428.950 ;
    RECT 0 429.410 0.460 429.410 ;
    RECT 0 429.870 0.460 429.870 ;
    RECT 0 430.330 0.460 430.330 ;
    RECT 0 430.790 0.460 430.790 ;
    RECT 0 431.250 0.460 431.250 ;
    RECT 0 431.710 0.460 431.710 ;
    RECT 0 432.170 0.460 432.170 ;
    RECT 0 432.630 0.460 432.630 ;
    RECT 0 433.090 0.460 433.090 ;
    RECT 0 433.550 0.460 433.550 ;
    RECT 0 434.010 0.460 434.010 ;
    RECT 0 434.470 0.460 434.470 ;
    RECT 0 434.930 0.460 434.930 ;
    RECT 0 435.390 0.460 435.390 ;
    RECT 0 435.850 0.460 435.850 ;
    RECT 0 436.310 0.460 436.310 ;
    RECT 0 436.770 0.460 436.770 ;
    RECT 0 437.230 0.460 437.230 ;
    RECT 0 437.690 0.460 437.690 ;
    RECT 0 438.150 0.460 438.150 ;
    RECT 0 438.610 0.460 438.610 ;
    RECT 0 439.070 0.460 439.070 ;
    RECT 0 439.530 0.460 439.530 ;
    RECT 0 439.990 0.460 439.990 ;
    RECT 0 440.450 0.460 440.450 ;
    RECT 0 440.910 0.460 440.910 ;
    RECT 0 441.370 0.460 441.370 ;
    RECT 0 441.830 0.460 441.830 ;
    RECT 0 442.290 0.460 442.290 ;
    RECT 0 442.750 0.460 442.750 ;
    RECT 0 443.210 0.460 443.210 ;
    RECT 0 443.670 0.460 443.670 ;
    RECT 0 444.130 0.460 444.130 ;
    RECT 0 444.590 0.460 444.590 ;
    RECT 0 445.050 0.460 445.050 ;
    RECT 0 445.510 0.460 445.510 ;
    RECT 0 445.970 0.460 445.970 ;
    RECT 0 446.430 0.460 446.430 ;
    RECT 0 446.890 0.460 446.890 ;
    RECT 0 447.350 0.460 447.350 ;
    RECT 0 447.810 0.460 447.810 ;
    RECT 0 448.270 0.460 448.270 ;
    RECT 0 448.730 0.460 448.730 ;
    RECT 0 449.190 0.460 449.190 ;
    RECT 0 449.650 0.460 449.650 ;
    RECT 0 450.110 0.460 450.110 ;
    RECT 0 450.570 0.460 450.570 ;
    RECT 0 451.030 0.460 451.030 ;
    RECT 0 451.490 0.460 451.490 ;
    RECT 0 451.950 0.460 451.950 ;
    RECT 0 452.410 0.460 452.410 ;
    RECT 0 452.870 0.460 452.870 ;
    RECT 0 453.330 0.460 453.330 ;
    RECT 0 453.790 0.460 453.790 ;
    RECT 0 454.250 0.460 454.250 ;
    RECT 0 454.710 0.460 454.710 ;
    RECT 0 455.170 0.460 455.170 ;
    RECT 0 455.630 0.460 455.630 ;
    RECT 0 456.090 0.460 456.090 ;
    RECT 0 456.550 0.460 456.550 ;
    RECT 0 457.010 0.460 457.010 ;
    RECT 0 457.470 0.460 457.470 ;
    RECT 0 457.930 0.460 457.930 ;
    RECT 0 458.390 0.460 458.390 ;
    RECT 0 458.850 0.460 458.850 ;
    RECT 0 459.310 0.460 459.310 ;
    RECT 0 459.770 0.460 459.770 ;
    RECT 0 460.230 0.460 460.230 ;
    RECT 0 460.690 0.460 460.690 ;
    RECT 0 461.150 0.460 461.150 ;
    RECT 0 461.610 0.460 461.610 ;
    RECT 0 462.070 0.460 462.070 ;
    RECT 0 462.530 0.460 462.530 ;
    RECT 0 462.990 0.460 462.990 ;
    RECT 0 463.450 0.460 463.450 ;
    RECT 0 463.910 0.460 463.910 ;
    RECT 0 464.370 0.460 464.370 ;
    RECT 0 464.830 0.460 464.830 ;
    RECT 0 465.290 0.460 465.290 ;
    RECT 0 465.750 0.460 465.750 ;
    RECT 0 466.210 0.460 466.210 ;
    RECT 0 466.670 0.460 466.670 ;
    RECT 0 467.130 0.460 467.130 ;
    RECT 0 467.590 0.460 467.590 ;
    RECT 0 468.050 0.460 468.050 ;
    RECT 0 468.510 0.460 468.510 ;
    RECT 0 468.970 0.460 468.970 ;
    RECT 0 469.430 0.460 469.430 ;
    RECT 0 469.890 0.460 469.890 ;
    RECT 0 470.350 0.460 470.350 ;
    RECT 0 470.810 0.460 470.810 ;
    RECT 0 471.270 0.460 471.270 ;
    RECT 0 471.730 0.460 471.730 ;
    RECT 0 472.190 0.460 472.190 ;
    RECT 0 472.650 0.460 472.650 ;
    RECT 0 473.110 0.460 473.110 ;
    RECT 0 473.570 0.460 473.570 ;
    RECT 0 474.030 0.460 474.030 ;
    RECT 0 474.490 0.460 474.490 ;
    RECT 0 474.950 0.460 474.950 ;
    RECT 0 475.410 0.460 475.410 ;
    RECT 0 475.870 0.460 475.870 ;
    RECT 0 476.330 0.460 476.330 ;
    RECT 0 476.790 0.460 476.790 ;
    RECT 0 477.250 0.460 477.250 ;
    RECT 0 477.710 0.460 477.710 ;
    RECT 0 478.170 0.460 478.170 ;
    RECT 0 478.630 0.460 478.630 ;
    RECT 0 479.090 0.460 479.090 ;
    RECT 0 479.550 0.460 479.550 ;
    RECT 0 480.010 0.460 480.010 ;
    RECT 0 480.470 0.460 480.470 ;
    RECT 0 480.930 0.460 480.930 ;
    RECT 0 481.390 0.460 481.390 ;
    RECT 0 481.850 0.460 481.850 ;
    RECT 0 482.310 0.460 482.310 ;
    RECT 0 482.770 0.460 482.770 ;
    RECT 0 483.230 0.460 483.230 ;
    RECT 0 483.690 0.460 483.690 ;
    RECT 0 484.150 0.460 484.150 ;
    RECT 0 484.610 0.460 484.610 ;
    RECT 0 485.070 0.460 485.070 ;
    RECT 0 485.530 0.460 485.530 ;
    RECT 0 485.990 0.460 485.990 ;
    RECT 0 486.450 0.460 486.450 ;
    RECT 0 486.910 0.460 486.910 ;
    RECT 0 487.370 0.460 487.370 ;
    RECT 0 487.830 0.460 487.830 ;
    RECT 0 488.290 0.460 488.290 ;
    RECT 0 488.750 0.460 488.750 ;
    RECT 0 489.210 0.460 489.210 ;
    RECT 0 489.670 0.460 489.670 ;
    RECT 0 490.130 0.460 490.130 ;
    RECT 0 490.590 0.460 490.590 ;
    RECT 0 491.050 0.460 491.050 ;
    RECT 0 491.510 0.460 491.510 ;
    RECT 0 491.970 0.460 491.970 ;
    RECT 0 492.430 0.460 492.430 ;
    RECT 0 492.890 0.460 492.890 ;
    RECT 0 493.350 0.460 493.350 ;
    RECT 0 493.810 0.460 493.810 ;
    RECT 0 494.270 0.460 494.270 ;
    RECT 0 494.730 0.460 494.730 ;
    RECT 0 495.190 0.460 495.190 ;
    RECT 0 495.650 0.460 495.650 ;
    RECT 0 496.110 0.460 496.110 ;
    RECT 0 496.570 0.460 496.570 ;
    RECT 0 497.030 0.460 497.030 ;
    RECT 0 497.490 0.460 497.490 ;
    RECT 0 497.950 0.460 497.950 ;
    RECT 0 498.410 0.460 498.410 ;
    RECT 0 498.870 0.460 498.870 ;
    RECT 0 499.330 0.460 499.330 ;
    RECT 0 499.790 0.460 499.790 ;
    RECT 0 500.250 0.460 500.250 ;
    RECT 0 500.710 0.460 500.710 ;
    RECT 0 501.170 0.460 501.170 ;
    RECT 0 501.630 0.460 501.630 ;
    RECT 0 502.090 0.460 502.090 ;
    RECT 0 502.550 0.460 502.550 ;
    RECT 0 503.010 0.460 503.010 ;
    RECT 0 503.470 0.460 503.470 ;
    RECT 0 503.930 0.460 503.930 ;
    RECT 0 504.390 0.460 504.390 ;
    RECT 0 504.850 0.460 504.850 ;
    RECT 0 505.310 0.460 505.310 ;
    RECT 0 505.770 0.460 505.770 ;
    RECT 0 506.230 0.460 506.230 ;
    RECT 0 506.690 0.460 506.690 ;
    RECT 0 507.150 0.460 507.150 ;
    RECT 0 507.610 0.460 507.610 ;
    RECT 0 508.070 0.460 508.070 ;
    RECT 0 508.530 0.460 508.530 ;
    RECT 0 508.990 0.460 508.990 ;
    RECT 0 509.450 0.460 509.450 ;
    RECT 0 509.910 0.460 509.910 ;
    RECT 0 510.370 0.460 510.370 ;
    RECT 0 510.830 0.460 510.830 ;
    RECT 0 511.290 0.460 511.290 ;
    RECT 0 511.750 0.460 511.750 ;
    RECT 0 512.210 0.460 512.210 ;
    RECT 0 512.670 0.460 512.670 ;
    RECT 0 513.130 0.460 513.130 ;
    RECT 0 513.590 0.460 513.590 ;
    RECT 0 514.050 0.460 514.050 ;
    RECT 0 514.510 0.460 514.510 ;
    RECT 0 514.970 0.460 514.970 ;
    RECT 0 515.430 0.460 515.430 ;
    RECT 0 515.890 0.460 515.890 ;
    RECT 0 516.350 0.460 516.350 ;
    RECT 0 516.810 0.460 516.810 ;
    RECT 0 517.270 0.460 517.270 ;
    RECT 0 517.730 0.460 517.730 ;
    RECT 0 518.190 0.460 518.190 ;
    RECT 0 518.650 0.460 518.650 ;
    RECT 0 519.110 0.460 519.110 ;
    RECT 0 519.570 0.460 519.570 ;
    RECT 0 520.030 0.460 520.030 ;
    RECT 0 520.490 0.460 520.490 ;
    RECT 0 520.950 0.460 520.950 ;
    RECT 0 521.410 0.460 521.410 ;
    RECT 0 521.870 0.460 521.870 ;
    RECT 0 522.330 0.460 522.330 ;
    RECT 0 522.790 0.460 522.790 ;
    RECT 0 523.250 0.460 523.250 ;
    RECT 0 523.710 0.460 523.710 ;
    RECT 0 524.170 0.460 524.170 ;
    RECT 0 524.630 0.460 524.630 ;
    RECT 0 525.090 0.460 525.090 ;
    RECT 0 525.550 0.460 525.550 ;
    RECT 0 526.010 0.460 526.010 ;
    RECT 0 526.470 0.460 526.470 ;
    RECT 0 526.930 0.460 526.930 ;
    RECT 0 527.390 0.460 527.390 ;
    RECT 0 527.850 0.460 527.850 ;
    RECT 0 528.310 0.460 528.310 ;
    RECT 0 528.770 0.460 528.770 ;
    RECT 0 529.230 0.460 529.230 ;
    RECT 0 529.690 0.460 529.690 ;
    RECT 0 530.150 0.460 530.150 ;
    RECT 0 530.610 0.460 530.610 ;
    RECT 0 531.070 0.460 531.070 ;
    RECT 0 531.530 0.460 531.530 ;
    RECT 0 531.990 0.460 531.990 ;
    RECT 0 532.450 0.460 532.450 ;
    RECT 0 532.910 0.460 532.910 ;
    RECT 0 533.370 0.460 533.370 ;
    RECT 0 533.830 0.460 533.830 ;
    RECT 0 534.290 0.460 534.290 ;
    RECT 0 534.750 0.460 534.750 ;
    RECT 0 535.210 0.460 535.210 ;
    RECT 0 535.670 0.460 535.670 ;
    RECT 0 536.130 0.460 536.130 ;
    RECT 0 536.590 0.460 536.590 ;
    RECT 0 537.050 0.460 537.050 ;
    RECT 0 537.510 0.460 537.510 ;
    RECT 0 537.970 0.460 537.970 ;
    RECT 0 538.430 0.460 538.430 ;
    RECT 0 538.890 0.460 538.890 ;
    RECT 0 539.350 0.460 539.350 ;
    RECT 0 539.810 0.460 539.810 ;
    RECT 0 540.270 0.460 540.270 ;
    RECT 0 540.730 0.460 540.730 ;
    RECT 0 541.190 0.460 541.190 ;
    RECT 0 541.650 0.460 541.650 ;
    RECT 0 542.110 0.460 542.110 ;
    RECT 0 542.570 0.460 542.570 ;
    RECT 0 543.030 0.460 543.030 ;
    RECT 0 543.490 0.460 543.490 ;
    RECT 0 543.950 0.460 543.950 ;
    RECT 0 544.410 0.460 544.410 ;
    RECT 0 544.870 0.460 544.870 ;
    RECT 0 545.330 0.460 545.330 ;
    RECT 0 545.790 0.460 545.790 ;
    RECT 0 546.250 0.460 546.250 ;
    RECT 0 546.710 0.460 546.710 ;
    RECT 0 547.170 0.460 547.170 ;
    RECT 0 547.630 0.460 547.630 ;
    RECT 0 548.090 0.460 548.090 ;
    RECT 0 548.550 0.460 548.550 ;
    RECT 0 549.010 0.460 549.010 ;
    RECT 0 549.470 0.460 549.470 ;
    RECT 0 549.930 0.460 549.930 ;
    RECT 0 550.390 0.460 550.390 ;
    RECT 0 550.850 0.460 550.850 ;
    RECT 0 551.310 0.460 551.310 ;
    RECT 0 551.770 0.460 551.770 ;
    RECT 0 552.230 0.460 552.230 ;
    RECT 0 552.690 0.460 552.690 ;
    RECT 0 553.150 0.460 553.150 ;
    RECT 0 553.610 0.460 553.610 ;
    RECT 0 554.070 0.460 554.070 ;
    RECT 0 554.530 0.460 554.530 ;
    RECT 0 554.990 0.460 554.990 ;
    RECT 0 555.450 0.460 555.450 ;
    RECT 0 555.910 0.460 555.910 ;
    RECT 0 556.370 0.460 556.370 ;
    RECT 0 556.830 0.460 556.830 ;
    RECT 0 557.290 0.460 557.290 ;
    RECT 0 557.750 0.460 640.090 ;
    RECT 0 640.550 0.460 640.550 ;
    RECT 0 641.010 0.460 641.010 ;
    RECT 0 641.470 0.460 641.470 ;
    RECT 0 641.930 0.460 641.930 ;
    RECT 0 642.390 0.460 642.390 ;
    RECT 0 642.850 0.460 642.850 ;
    RECT 0 643.310 0.460 643.310 ;
    RECT 0 643.770 0.460 643.770 ;
    RECT 0 644.230 0.460 644.230 ;
    RECT 0 644.690 0.460 644.690 ;
    RECT 0 645.150 0.460 645.150 ;
    RECT 0 645.610 0.460 645.610 ;
    RECT 0 646.070 0.460 646.070 ;
    RECT 0 646.530 0.460 646.530 ;
    RECT 0 646.990 0.460 646.990 ;
    RECT 0 647.450 0.460 647.450 ;
    RECT 0 647.910 0.460 647.910 ;
    RECT 0 648.370 0.460 648.370 ;
    RECT 0 648.830 0.460 648.830 ;
    RECT 0 649.290 0.460 649.290 ;
    RECT 0 649.750 0.460 649.750 ;
    RECT 0 650.210 0.460 650.210 ;
    RECT 0 650.670 0.460 650.670 ;
    RECT 0 651.130 0.460 651.130 ;
    RECT 0 651.590 0.460 651.590 ;
    RECT 0 652.050 0.460 652.050 ;
    RECT 0 652.510 0.460 652.510 ;
    RECT 0 652.970 0.460 652.970 ;
    RECT 0 653.430 0.460 653.430 ;
    RECT 0 653.890 0.460 653.890 ;
    RECT 0 654.350 0.460 654.350 ;
    RECT 0 654.810 0.460 654.810 ;
    RECT 0 655.270 0.460 655.270 ;
    RECT 0 655.730 0.460 655.730 ;
    RECT 0 656.190 0.460 656.190 ;
    RECT 0 656.650 0.460 656.650 ;
    RECT 0 657.110 0.460 657.110 ;
    RECT 0 657.570 0.460 657.570 ;
    RECT 0 658.030 0.460 658.030 ;
    RECT 0 658.490 0.460 658.490 ;
    RECT 0 658.950 0.460 658.950 ;
    RECT 0 659.410 0.460 659.410 ;
    RECT 0 659.870 0.460 659.870 ;
    RECT 0 660.330 0.460 660.330 ;
    RECT 0 660.790 0.460 660.790 ;
    RECT 0 661.250 0.460 661.250 ;
    RECT 0 661.710 0.460 661.710 ;
    RECT 0 662.170 0.460 662.170 ;
    RECT 0 662.630 0.460 662.630 ;
    RECT 0 663.090 0.460 663.090 ;
    RECT 0 663.550 0.460 663.550 ;
    RECT 0 664.010 0.460 664.010 ;
    RECT 0 664.470 0.460 664.470 ;
    RECT 0 664.930 0.460 664.930 ;
    RECT 0 665.390 0.460 665.390 ;
    RECT 0 665.850 0.460 665.850 ;
    RECT 0 666.310 0.460 666.310 ;
    RECT 0 666.770 0.460 666.770 ;
    RECT 0 667.230 0.460 667.230 ;
    RECT 0 667.690 0.460 667.690 ;
    RECT 0 668.150 0.460 668.150 ;
    RECT 0 668.610 0.460 668.610 ;
    RECT 0 669.070 0.460 669.070 ;
    RECT 0 669.530 0.460 669.530 ;
    RECT 0 669.990 0.460 669.990 ;
    RECT 0 670.450 0.460 670.450 ;
    RECT 0 670.910 0.460 670.910 ;
    RECT 0 671.370 0.460 671.370 ;
    RECT 0 671.830 0.460 671.830 ;
    RECT 0 672.290 0.460 672.290 ;
    RECT 0 672.750 0.460 672.750 ;
    RECT 0 673.210 0.460 673.210 ;
    RECT 0 673.670 0.460 673.670 ;
    RECT 0 674.130 0.460 674.130 ;
    RECT 0 674.590 0.460 674.590 ;
    RECT 0 675.050 0.460 675.050 ;
    RECT 0 675.510 0.460 675.510 ;
    RECT 0 675.970 0.460 675.970 ;
    RECT 0 676.430 0.460 676.430 ;
    RECT 0 676.890 0.460 676.890 ;
    RECT 0 677.350 0.460 677.350 ;
    RECT 0 677.810 0.460 677.810 ;
    RECT 0 678.270 0.460 678.270 ;
    RECT 0 678.730 0.460 678.730 ;
    RECT 0 679.190 0.460 679.190 ;
    RECT 0 679.650 0.460 679.650 ;
    RECT 0 680.110 0.460 680.110 ;
    RECT 0 680.570 0.460 680.570 ;
    RECT 0 681.030 0.460 681.030 ;
    RECT 0 681.490 0.460 681.490 ;
    RECT 0 681.950 0.460 681.950 ;
    RECT 0 682.410 0.460 682.410 ;
    RECT 0 682.870 0.460 682.870 ;
    RECT 0 683.330 0.460 683.330 ;
    RECT 0 683.790 0.460 683.790 ;
    RECT 0 684.250 0.460 684.250 ;
    RECT 0 684.710 0.460 684.710 ;
    RECT 0 685.170 0.460 685.170 ;
    RECT 0 685.630 0.460 685.630 ;
    RECT 0 686.090 0.460 686.090 ;
    RECT 0 686.550 0.460 686.550 ;
    RECT 0 687.010 0.460 687.010 ;
    RECT 0 687.470 0.460 687.470 ;
    RECT 0 687.930 0.460 687.930 ;
    RECT 0 688.390 0.460 688.390 ;
    RECT 0 688.850 0.460 688.850 ;
    RECT 0 689.310 0.460 689.310 ;
    RECT 0 689.770 0.460 689.770 ;
    RECT 0 690.230 0.460 690.230 ;
    RECT 0 690.690 0.460 690.690 ;
    RECT 0 691.150 0.460 691.150 ;
    RECT 0 691.610 0.460 691.610 ;
    RECT 0 692.070 0.460 692.070 ;
    RECT 0 692.530 0.460 692.530 ;
    RECT 0 692.990 0.460 692.990 ;
    RECT 0 693.450 0.460 693.450 ;
    RECT 0 693.910 0.460 693.910 ;
    RECT 0 694.370 0.460 694.370 ;
    RECT 0 694.830 0.460 694.830 ;
    RECT 0 695.290 0.460 695.290 ;
    RECT 0 695.750 0.460 695.750 ;
    RECT 0 696.210 0.460 696.210 ;
    RECT 0 696.670 0.460 696.670 ;
    RECT 0 697.130 0.460 697.130 ;
    RECT 0 697.590 0.460 697.590 ;
    RECT 0 698.050 0.460 698.050 ;
    RECT 0 698.510 0.460 698.510 ;
    RECT 0 698.970 0.460 698.970 ;
    RECT 0 699.430 0.460 699.430 ;
    RECT 0 699.890 0.460 699.890 ;
    RECT 0 700.350 0.460 700.350 ;
    RECT 0 700.810 0.460 700.810 ;
    RECT 0 701.270 0.460 701.270 ;
    RECT 0 701.730 0.460 701.730 ;
    RECT 0 702.190 0.460 702.190 ;
    RECT 0 702.650 0.460 702.650 ;
    RECT 0 703.110 0.460 703.110 ;
    RECT 0 703.570 0.460 703.570 ;
    RECT 0 704.030 0.460 704.030 ;
    RECT 0 704.490 0.460 704.490 ;
    RECT 0 704.950 0.460 704.950 ;
    RECT 0 705.410 0.460 705.410 ;
    RECT 0 705.870 0.460 705.870 ;
    RECT 0 706.330 0.460 706.330 ;
    RECT 0 706.790 0.460 706.790 ;
    RECT 0 707.250 0.460 707.250 ;
    RECT 0 707.710 0.460 707.710 ;
    RECT 0 708.170 0.460 708.170 ;
    RECT 0 708.630 0.460 708.630 ;
    RECT 0 709.090 0.460 709.090 ;
    RECT 0 709.550 0.460 709.550 ;
    RECT 0 710.010 0.460 710.010 ;
    RECT 0 710.470 0.460 710.470 ;
    RECT 0 710.930 0.460 710.930 ;
    RECT 0 711.390 0.460 711.390 ;
    RECT 0 711.850 0.460 711.850 ;
    RECT 0 712.310 0.460 712.310 ;
    RECT 0 712.770 0.460 712.770 ;
    RECT 0 713.230 0.460 713.230 ;
    RECT 0 713.690 0.460 713.690 ;
    RECT 0 714.150 0.460 714.150 ;
    RECT 0 714.610 0.460 714.610 ;
    RECT 0 715.070 0.460 715.070 ;
    RECT 0 715.530 0.460 715.530 ;
    RECT 0 715.990 0.460 715.990 ;
    RECT 0 716.450 0.460 716.450 ;
    RECT 0 716.910 0.460 716.910 ;
    RECT 0 717.370 0.460 717.370 ;
    RECT 0 717.830 0.460 717.830 ;
    RECT 0 718.290 0.460 718.290 ;
    RECT 0 718.750 0.460 718.750 ;
    RECT 0 719.210 0.460 719.210 ;
    RECT 0 719.670 0.460 719.670 ;
    RECT 0 720.130 0.460 720.130 ;
    RECT 0 720.590 0.460 720.590 ;
    RECT 0 721.050 0.460 721.050 ;
    RECT 0 721.510 0.460 721.510 ;
    RECT 0 721.970 0.460 721.970 ;
    RECT 0 722.430 0.460 722.430 ;
    RECT 0 722.890 0.460 722.890 ;
    RECT 0 723.350 0.460 723.350 ;
    RECT 0 723.810 0.460 723.810 ;
    RECT 0 724.270 0.460 724.270 ;
    RECT 0 724.730 0.460 724.730 ;
    RECT 0 725.190 0.460 725.190 ;
    RECT 0 725.650 0.460 725.650 ;
    RECT 0 726.110 0.460 726.110 ;
    RECT 0 726.570 0.460 726.570 ;
    RECT 0 727.030 0.460 727.030 ;
    RECT 0 727.490 0.460 727.490 ;
    RECT 0 727.950 0.460 727.950 ;
    RECT 0 728.410 0.460 728.410 ;
    RECT 0 728.870 0.460 728.870 ;
    RECT 0 729.330 0.460 729.330 ;
    RECT 0 729.790 0.460 729.790 ;
    RECT 0 730.250 0.460 730.250 ;
    RECT 0 730.710 0.460 730.710 ;
    RECT 0 731.170 0.460 731.170 ;
    RECT 0 731.630 0.460 731.630 ;
    RECT 0 732.090 0.460 732.090 ;
    RECT 0 732.550 0.460 732.550 ;
    RECT 0 733.010 0.460 733.010 ;
    RECT 0 733.470 0.460 733.470 ;
    RECT 0 733.930 0.460 733.930 ;
    RECT 0 734.390 0.460 734.390 ;
    RECT 0 734.850 0.460 734.850 ;
    RECT 0 735.310 0.460 735.310 ;
    RECT 0 735.770 0.460 735.770 ;
    RECT 0 736.230 0.460 736.230 ;
    RECT 0 736.690 0.460 736.690 ;
    RECT 0 737.150 0.460 737.150 ;
    RECT 0 737.610 0.460 737.610 ;
    RECT 0 738.070 0.460 738.070 ;
    RECT 0 738.530 0.460 738.530 ;
    RECT 0 738.990 0.460 738.990 ;
    RECT 0 739.450 0.460 739.450 ;
    RECT 0 739.910 0.460 739.910 ;
    RECT 0 740.370 0.460 740.370 ;
    RECT 0 740.830 0.460 740.830 ;
    RECT 0 741.290 0.460 741.290 ;
    RECT 0 741.750 0.460 741.750 ;
    RECT 0 742.210 0.460 742.210 ;
    RECT 0 742.670 0.460 742.670 ;
    RECT 0 743.130 0.460 743.130 ;
    RECT 0 743.590 0.460 743.590 ;
    RECT 0 744.050 0.460 744.050 ;
    RECT 0 744.510 0.460 744.510 ;
    RECT 0 744.970 0.460 744.970 ;
    RECT 0 745.430 0.460 745.430 ;
    RECT 0 745.890 0.460 745.890 ;
    RECT 0 746.350 0.460 746.350 ;
    RECT 0 746.810 0.460 746.810 ;
    RECT 0 747.270 0.460 747.270 ;
    RECT 0 747.730 0.460 747.730 ;
    RECT 0 748.190 0.460 748.190 ;
    RECT 0 748.650 0.460 748.650 ;
    RECT 0 749.110 0.460 749.110 ;
    RECT 0 749.570 0.460 749.570 ;
    RECT 0 750.030 0.460 750.030 ;
    RECT 0 750.490 0.460 750.490 ;
    RECT 0 750.950 0.460 750.950 ;
    RECT 0 751.410 0.460 751.410 ;
    RECT 0 751.870 0.460 751.870 ;
    RECT 0 752.330 0.460 752.330 ;
    RECT 0 752.790 0.460 752.790 ;
    RECT 0 753.250 0.460 753.250 ;
    RECT 0 753.710 0.460 753.710 ;
    RECT 0 754.170 0.460 754.170 ;
    RECT 0 754.630 0.460 754.630 ;
    RECT 0 755.090 0.460 755.090 ;
    RECT 0 755.550 0.460 755.550 ;
    RECT 0 756.010 0.460 756.010 ;
    RECT 0 756.470 0.460 756.470 ;
    RECT 0 756.930 0.460 756.930 ;
    RECT 0 757.390 0.460 757.390 ;
    RECT 0 757.850 0.460 757.850 ;
    RECT 0 758.310 0.460 758.310 ;
    RECT 0 758.770 0.460 758.770 ;
    RECT 0 759.230 0.460 759.230 ;
    RECT 0 759.690 0.460 759.690 ;
    RECT 0 760.150 0.460 760.150 ;
    RECT 0 760.610 0.460 760.610 ;
    RECT 0 761.070 0.460 761.070 ;
    RECT 0 761.530 0.460 761.530 ;
    RECT 0 761.990 0.460 761.990 ;
    RECT 0 762.450 0.460 762.450 ;
    RECT 0 762.910 0.460 762.910 ;
    RECT 0 763.370 0.460 763.370 ;
    RECT 0 763.830 0.460 763.830 ;
    RECT 0 764.290 0.460 764.290 ;
    RECT 0 764.750 0.460 764.750 ;
    RECT 0 765.210 0.460 765.210 ;
    RECT 0 765.670 0.460 765.670 ;
    RECT 0 766.130 0.460 766.130 ;
    RECT 0 766.590 0.460 766.590 ;
    RECT 0 767.050 0.460 767.050 ;
    RECT 0 767.510 0.460 767.510 ;
    RECT 0 767.970 0.460 767.970 ;
    RECT 0 768.430 0.460 768.430 ;
    RECT 0 768.890 0.460 768.890 ;
    RECT 0 769.350 0.460 769.350 ;
    RECT 0 769.810 0.460 769.810 ;
    RECT 0 770.270 0.460 770.270 ;
    RECT 0 770.730 0.460 770.730 ;
    RECT 0 771.190 0.460 771.190 ;
    RECT 0 771.650 0.460 771.650 ;
    RECT 0 772.110 0.460 772.110 ;
    RECT 0 772.570 0.460 772.570 ;
    RECT 0 773.030 0.460 773.030 ;
    RECT 0 773.490 0.460 773.490 ;
    RECT 0 773.950 0.460 773.950 ;
    RECT 0 774.410 0.460 774.410 ;
    RECT 0 774.870 0.460 774.870 ;
    RECT 0 775.330 0.460 775.330 ;
    RECT 0 775.790 0.460 775.790 ;
    RECT 0 776.250 0.460 776.250 ;
    RECT 0 776.710 0.460 776.710 ;
    RECT 0 777.170 0.460 777.170 ;
    RECT 0 777.630 0.460 777.630 ;
    RECT 0 778.090 0.460 778.090 ;
    RECT 0 778.550 0.460 778.550 ;
    RECT 0 779.010 0.460 779.010 ;
    RECT 0 779.470 0.460 779.470 ;
    RECT 0 779.930 0.460 779.930 ;
    RECT 0 780.390 0.460 780.390 ;
    RECT 0 780.850 0.460 780.850 ;
    RECT 0 781.310 0.460 781.310 ;
    RECT 0 781.770 0.460 781.770 ;
    RECT 0 782.230 0.460 782.230 ;
    RECT 0 782.690 0.460 782.690 ;
    RECT 0 783.150 0.460 783.150 ;
    RECT 0 783.610 0.460 783.610 ;
    RECT 0 784.070 0.460 784.070 ;
    RECT 0 784.530 0.460 784.530 ;
    RECT 0 784.990 0.460 784.990 ;
    RECT 0 785.450 0.460 785.450 ;
    RECT 0 785.910 0.460 785.910 ;
    RECT 0 786.370 0.460 786.370 ;
    RECT 0 786.830 0.460 786.830 ;
    RECT 0 787.290 0.460 787.290 ;
    RECT 0 787.750 0.460 787.750 ;
    RECT 0 788.210 0.460 788.210 ;
    RECT 0 788.670 0.460 788.670 ;
    RECT 0 789.130 0.460 789.130 ;
    RECT 0 789.590 0.460 789.590 ;
    RECT 0 790.050 0.460 790.050 ;
    RECT 0 790.510 0.460 790.510 ;
    RECT 0 790.970 0.460 790.970 ;
    RECT 0 791.430 0.460 791.430 ;
    RECT 0 791.890 0.460 791.890 ;
    RECT 0 792.350 0.460 792.350 ;
    RECT 0 792.810 0.460 792.810 ;
    RECT 0 793.270 0.460 793.270 ;
    RECT 0 793.730 0.460 793.730 ;
    RECT 0 794.190 0.460 794.190 ;
    RECT 0 794.650 0.460 794.650 ;
    RECT 0 795.110 0.460 795.110 ;
    RECT 0 795.570 0.460 795.570 ;
    RECT 0 796.030 0.460 796.030 ;
    RECT 0 796.490 0.460 796.490 ;
    RECT 0 796.950 0.460 796.950 ;
    RECT 0 797.410 0.460 797.410 ;
    RECT 0 797.870 0.460 797.870 ;
    RECT 0 798.330 0.460 798.330 ;
    RECT 0 798.790 0.460 798.790 ;
    RECT 0 799.250 0.460 799.250 ;
    RECT 0 799.710 0.460 799.710 ;
    RECT 0 800.170 0.460 800.170 ;
    RECT 0 800.630 0.460 800.630 ;
    RECT 0 801.090 0.460 801.090 ;
    RECT 0 801.550 0.460 801.550 ;
    RECT 0 802.010 0.460 802.010 ;
    RECT 0 802.470 0.460 802.470 ;
    RECT 0 802.930 0.460 802.930 ;
    RECT 0 803.390 0.460 803.390 ;
    RECT 0 803.850 0.460 803.850 ;
    RECT 0 804.310 0.460 804.310 ;
    RECT 0 804.770 0.460 804.770 ;
    RECT 0 805.230 0.460 805.230 ;
    RECT 0 805.690 0.460 805.690 ;
    RECT 0 806.150 0.460 806.150 ;
    RECT 0 806.610 0.460 806.610 ;
    RECT 0 807.070 0.460 807.070 ;
    RECT 0 807.530 0.460 807.530 ;
    RECT 0 807.990 0.460 807.990 ;
    RECT 0 808.450 0.460 808.450 ;
    RECT 0 808.910 0.460 808.910 ;
    RECT 0 809.370 0.460 809.370 ;
    RECT 0 809.830 0.460 809.830 ;
    RECT 0 810.290 0.460 810.290 ;
    RECT 0 810.750 0.460 810.750 ;
    RECT 0 811.210 0.460 811.210 ;
    RECT 0 811.670 0.460 811.670 ;
    RECT 0 812.130 0.460 812.130 ;
    RECT 0 812.590 0.460 812.590 ;
    RECT 0 813.050 0.460 813.050 ;
    RECT 0 813.510 0.460 813.510 ;
    RECT 0 813.970 0.460 813.970 ;
    RECT 0 814.430 0.460 814.430 ;
    RECT 0 814.890 0.460 814.890 ;
    RECT 0 815.350 0.460 815.350 ;
    RECT 0 815.810 0.460 815.810 ;
    RECT 0 816.270 0.460 816.270 ;
    RECT 0 816.730 0.460 816.730 ;
    RECT 0 817.190 0.460 817.190 ;
    RECT 0 817.650 0.460 817.650 ;
    RECT 0 818.110 0.460 818.110 ;
    RECT 0 818.570 0.460 818.570 ;
    RECT 0 819.030 0.460 819.030 ;
    RECT 0 819.490 0.460 819.490 ;
    RECT 0 819.950 0.460 819.950 ;
    RECT 0 820.410 0.460 820.410 ;
    RECT 0 820.870 0.460 820.870 ;
    RECT 0 821.330 0.460 821.330 ;
    RECT 0 821.790 0.460 821.790 ;
    RECT 0 822.250 0.460 822.250 ;
    RECT 0 822.710 0.460 822.710 ;
    RECT 0 823.170 0.460 823.170 ;
    RECT 0 823.630 0.460 823.630 ;
    RECT 0 824.090 0.460 824.090 ;
    RECT 0 824.550 0.460 824.550 ;
    RECT 0 825.010 0.460 825.010 ;
    RECT 0 825.470 0.460 825.470 ;
    RECT 0 825.930 0.460 825.930 ;
    RECT 0 826.390 0.460 826.390 ;
    RECT 0 826.850 0.460 826.850 ;
    RECT 0 827.310 0.460 827.310 ;
    RECT 0 827.770 0.460 827.770 ;
    RECT 0 828.230 0.460 828.230 ;
    RECT 0 828.690 0.460 828.690 ;
    RECT 0 829.150 0.460 829.150 ;
    RECT 0 829.610 0.460 829.610 ;
    RECT 0 830.070 0.460 830.070 ;
    RECT 0 830.530 0.460 830.530 ;
    RECT 0 830.990 0.460 830.990 ;
    RECT 0 831.450 0.460 831.450 ;
    RECT 0 831.910 0.460 831.910 ;
    RECT 0 832.370 0.460 832.370 ;
    RECT 0 832.830 0.460 832.830 ;
    RECT 0 833.290 0.460 833.290 ;
    RECT 0 833.750 0.460 833.750 ;
    RECT 0 834.210 0.460 834.210 ;
    RECT 0 834.670 0.460 834.670 ;
    RECT 0 835.130 0.460 835.130 ;
    RECT 0 835.590 0.460 835.590 ;
    RECT 0 836.050 0.460 836.050 ;
    RECT 0 836.510 0.460 836.510 ;
    RECT 0 836.970 0.460 836.970 ;
    RECT 0 837.430 0.460 837.430 ;
    RECT 0 837.890 0.460 837.890 ;
    RECT 0 838.350 0.460 838.350 ;
    RECT 0 838.810 0.460 838.810 ;
    RECT 0 839.270 0.460 839.270 ;
    RECT 0 839.730 0.460 839.730 ;
    RECT 0 840.190 0.460 840.190 ;
    RECT 0 840.650 0.460 840.650 ;
    RECT 0 841.110 0.460 841.110 ;
    RECT 0 841.570 0.460 841.570 ;
    RECT 0 842.030 0.460 842.030 ;
    RECT 0 842.490 0.460 842.490 ;
    RECT 0 842.950 0.460 842.950 ;
    RECT 0 843.410 0.460 843.410 ;
    RECT 0 843.870 0.460 843.870 ;
    RECT 0 844.330 0.460 844.330 ;
    RECT 0 844.790 0.460 844.790 ;
    RECT 0 845.250 0.460 845.250 ;
    RECT 0 845.710 0.460 845.710 ;
    RECT 0 846.170 0.460 846.170 ;
    RECT 0 846.630 0.460 846.630 ;
    RECT 0 847.090 0.460 847.090 ;
    RECT 0 847.550 0.460 847.550 ;
    RECT 0 848.010 0.460 848.010 ;
    RECT 0 848.470 0.460 848.470 ;
    RECT 0 848.930 0.460 848.930 ;
    RECT 0 849.390 0.460 849.390 ;
    RECT 0 849.850 0.460 849.850 ;
    RECT 0 850.310 0.460 850.310 ;
    RECT 0 850.770 0.460 850.770 ;
    RECT 0 851.230 0.460 851.230 ;
    RECT 0 851.690 0.460 851.690 ;
    RECT 0 852.150 0.460 852.150 ;
    RECT 0 852.610 0.460 852.610 ;
    RECT 0 853.070 0.460 853.070 ;
    RECT 0 853.530 0.460 853.530 ;
    RECT 0 853.990 0.460 853.990 ;
    RECT 0 854.450 0.460 854.450 ;
    RECT 0 854.910 0.460 854.910 ;
    RECT 0 855.370 0.460 855.370 ;
    RECT 0 855.830 0.460 855.830 ;
    RECT 0 856.290 0.460 856.290 ;
    RECT 0 856.750 0.460 856.750 ;
    RECT 0 857.210 0.460 857.210 ;
    RECT 0 857.670 0.460 857.670 ;
    RECT 0 858.130 0.460 858.130 ;
    RECT 0 858.590 0.460 858.590 ;
    RECT 0 859.050 0.460 859.050 ;
    RECT 0 859.510 0.460 859.510 ;
    RECT 0 859.970 0.460 859.970 ;
    RECT 0 860.430 0.460 860.430 ;
    RECT 0 860.890 0.460 860.890 ;
    RECT 0 861.350 0.460 861.350 ;
    RECT 0 861.810 0.460 861.810 ;
    RECT 0 862.270 0.460 862.270 ;
    RECT 0 862.730 0.460 862.730 ;
    RECT 0 863.190 0.460 863.190 ;
    RECT 0 863.650 0.460 863.650 ;
    RECT 0 864.110 0.460 864.110 ;
    RECT 0 864.570 0.460 864.570 ;
    RECT 0 865.030 0.460 865.030 ;
    RECT 0 865.490 0.460 865.490 ;
    RECT 0 865.950 0.460 865.950 ;
    RECT 0 866.410 0.460 866.410 ;
    RECT 0 866.870 0.460 866.870 ;
    RECT 0 867.330 0.460 867.330 ;
    RECT 0 867.790 0.460 867.790 ;
    RECT 0 868.250 0.460 868.250 ;
    RECT 0 868.710 0.460 868.710 ;
    RECT 0 869.170 0.460 869.170 ;
    RECT 0 869.630 0.460 869.630 ;
    RECT 0 870.090 0.460 870.090 ;
    RECT 0 870.550 0.460 870.550 ;
    RECT 0 871.010 0.460 871.010 ;
    RECT 0 871.470 0.460 871.470 ;
    RECT 0 871.930 0.460 871.930 ;
    RECT 0 872.390 0.460 872.390 ;
    RECT 0 872.850 0.460 872.850 ;
    RECT 0 873.310 0.460 873.310 ;
    RECT 0 873.770 0.460 873.770 ;
    RECT 0 874.230 0.460 874.230 ;
    RECT 0 874.690 0.460 874.690 ;
    RECT 0 875.150 0.460 875.150 ;
    RECT 0 875.610 0.460 957.950 ;
    RECT 0 958.410 0.460 958.410 ;
    RECT 0 958.870 0.460 958.870 ;
    RECT 0 959.330 0.460 959.330 ;
    RECT 0 959.790 0.460 959.790 ;
    RECT 0 960.250 0.460 960.250 ;
    RECT 0 960.710 0.460 960.710 ;
    RECT 0 961.170 0.460 961.170 ;
    RECT 0 961.630 0.460 1043.970 ;
    RECT 0 1044.430 0.460 1044.430 ;
    RECT 0 1044.890 0.460 1044.890 ;
    RECT 0 1045.350 0.460 1052.640 ;
    LAYER met4 ;
    RECT 0 0 834.440 4.600 ;
    RECT 0 1048.040 834.440 1052.640 ;
    RECT 0.000 4.600 3.680 1048.040 ;
    RECT 5.520 4.600 7.360 1048.040 ;
    RECT 9.200 4.600 11.040 1048.040 ;
    RECT 12.880 4.600 14.720 1048.040 ;
    RECT 16.560 4.600 18.400 1048.040 ;
    RECT 20.240 4.600 22.080 1048.040 ;
    RECT 23.920 4.600 25.760 1048.040 ;
    RECT 27.600 4.600 29.440 1048.040 ;
    RECT 31.280 4.600 33.120 1048.040 ;
    RECT 34.960 4.600 36.800 1048.040 ;
    RECT 38.640 4.600 40.480 1048.040 ;
    RECT 42.320 4.600 44.160 1048.040 ;
    RECT 46.000 4.600 47.840 1048.040 ;
    RECT 49.680 4.600 51.520 1048.040 ;
    RECT 53.360 4.600 55.200 1048.040 ;
    RECT 57.040 4.600 58.880 1048.040 ;
    RECT 60.720 4.600 62.560 1048.040 ;
    RECT 64.400 4.600 66.240 1048.040 ;
    RECT 68.080 4.600 69.920 1048.040 ;
    RECT 71.760 4.600 73.600 1048.040 ;
    RECT 75.440 4.600 77.280 1048.040 ;
    RECT 79.120 4.600 80.960 1048.040 ;
    RECT 82.800 4.600 84.640 1048.040 ;
    RECT 86.480 4.600 88.320 1048.040 ;
    RECT 90.160 4.600 92.000 1048.040 ;
    RECT 93.840 4.600 95.680 1048.040 ;
    RECT 97.520 4.600 99.360 1048.040 ;
    RECT 101.200 4.600 103.040 1048.040 ;
    RECT 104.880 4.600 106.720 1048.040 ;
    RECT 108.560 4.600 110.400 1048.040 ;
    RECT 112.240 4.600 114.080 1048.040 ;
    RECT 115.920 4.600 117.760 1048.040 ;
    RECT 119.600 4.600 121.440 1048.040 ;
    RECT 123.280 4.600 125.120 1048.040 ;
    RECT 126.960 4.600 128.800 1048.040 ;
    RECT 130.640 4.600 132.480 1048.040 ;
    RECT 134.320 4.600 136.160 1048.040 ;
    RECT 138.000 4.600 139.840 1048.040 ;
    RECT 141.680 4.600 143.520 1048.040 ;
    RECT 145.360 4.600 147.200 1048.040 ;
    RECT 149.040 4.600 150.880 1048.040 ;
    RECT 152.720 4.600 154.560 1048.040 ;
    RECT 156.400 4.600 158.240 1048.040 ;
    RECT 160.080 4.600 161.920 1048.040 ;
    RECT 163.760 4.600 165.600 1048.040 ;
    RECT 167.440 4.600 169.280 1048.040 ;
    RECT 171.120 4.600 172.960 1048.040 ;
    RECT 174.800 4.600 176.640 1048.040 ;
    RECT 178.480 4.600 180.320 1048.040 ;
    RECT 182.160 4.600 184.000 1048.040 ;
    RECT 185.840 4.600 187.680 1048.040 ;
    RECT 189.520 4.600 191.360 1048.040 ;
    RECT 193.200 4.600 195.040 1048.040 ;
    RECT 196.880 4.600 198.720 1048.040 ;
    RECT 200.560 4.600 202.400 1048.040 ;
    RECT 204.240 4.600 206.080 1048.040 ;
    RECT 207.920 4.600 209.760 1048.040 ;
    RECT 211.600 4.600 213.440 1048.040 ;
    RECT 215.280 4.600 217.120 1048.040 ;
    RECT 218.960 4.600 220.800 1048.040 ;
    RECT 222.640 4.600 224.480 1048.040 ;
    RECT 226.320 4.600 228.160 1048.040 ;
    RECT 230.000 4.600 231.840 1048.040 ;
    RECT 233.680 4.600 235.520 1048.040 ;
    RECT 237.360 4.600 239.200 1048.040 ;
    RECT 241.040 4.600 242.880 1048.040 ;
    RECT 244.720 4.600 246.560 1048.040 ;
    RECT 248.400 4.600 250.240 1048.040 ;
    RECT 252.080 4.600 253.920 1048.040 ;
    RECT 255.760 4.600 257.600 1048.040 ;
    RECT 259.440 4.600 261.280 1048.040 ;
    RECT 263.120 4.600 264.960 1048.040 ;
    RECT 266.800 4.600 268.640 1048.040 ;
    RECT 270.480 4.600 272.320 1048.040 ;
    RECT 274.160 4.600 276.000 1048.040 ;
    RECT 277.840 4.600 279.680 1048.040 ;
    RECT 281.520 4.600 283.360 1048.040 ;
    RECT 285.200 4.600 287.040 1048.040 ;
    RECT 288.880 4.600 290.720 1048.040 ;
    RECT 292.560 4.600 294.400 1048.040 ;
    RECT 296.240 4.600 298.080 1048.040 ;
    RECT 299.920 4.600 301.760 1048.040 ;
    RECT 303.600 4.600 305.440 1048.040 ;
    RECT 307.280 4.600 309.120 1048.040 ;
    RECT 310.960 4.600 312.800 1048.040 ;
    RECT 314.640 4.600 316.480 1048.040 ;
    RECT 318.320 4.600 320.160 1048.040 ;
    RECT 322.000 4.600 323.840 1048.040 ;
    RECT 325.680 4.600 327.520 1048.040 ;
    RECT 329.360 4.600 331.200 1048.040 ;
    RECT 333.040 4.600 334.880 1048.040 ;
    RECT 336.720 4.600 338.560 1048.040 ;
    RECT 340.400 4.600 342.240 1048.040 ;
    RECT 344.080 4.600 345.920 1048.040 ;
    RECT 347.760 4.600 349.600 1048.040 ;
    RECT 351.440 4.600 353.280 1048.040 ;
    RECT 355.120 4.600 356.960 1048.040 ;
    RECT 358.800 4.600 360.640 1048.040 ;
    RECT 362.480 4.600 364.320 1048.040 ;
    RECT 366.160 4.600 368.000 1048.040 ;
    RECT 369.840 4.600 371.680 1048.040 ;
    RECT 373.520 4.600 375.360 1048.040 ;
    RECT 377.200 4.600 379.040 1048.040 ;
    RECT 380.880 4.600 382.720 1048.040 ;
    RECT 384.560 4.600 386.400 1048.040 ;
    RECT 388.240 4.600 390.080 1048.040 ;
    RECT 391.920 4.600 393.760 1048.040 ;
    RECT 395.600 4.600 397.440 1048.040 ;
    RECT 399.280 4.600 401.120 1048.040 ;
    RECT 402.960 4.600 404.800 1048.040 ;
    RECT 406.640 4.600 408.480 1048.040 ;
    RECT 410.320 4.600 412.160 1048.040 ;
    RECT 414.000 4.600 415.840 1048.040 ;
    RECT 417.680 4.600 419.520 1048.040 ;
    RECT 421.360 4.600 423.200 1048.040 ;
    RECT 425.040 4.600 426.880 1048.040 ;
    RECT 428.720 4.600 430.560 1048.040 ;
    RECT 432.400 4.600 434.240 1048.040 ;
    RECT 436.080 4.600 437.920 1048.040 ;
    RECT 439.760 4.600 441.600 1048.040 ;
    RECT 443.440 4.600 445.280 1048.040 ;
    RECT 447.120 4.600 448.960 1048.040 ;
    RECT 450.800 4.600 452.640 1048.040 ;
    RECT 454.480 4.600 456.320 1048.040 ;
    RECT 458.160 4.600 460.000 1048.040 ;
    RECT 461.840 4.600 463.680 1048.040 ;
    RECT 465.520 4.600 467.360 1048.040 ;
    RECT 469.200 4.600 471.040 1048.040 ;
    RECT 472.880 4.600 474.720 1048.040 ;
    RECT 476.560 4.600 478.400 1048.040 ;
    RECT 480.240 4.600 482.080 1048.040 ;
    RECT 483.920 4.600 485.760 1048.040 ;
    RECT 487.600 4.600 489.440 1048.040 ;
    RECT 491.280 4.600 493.120 1048.040 ;
    RECT 494.960 4.600 496.800 1048.040 ;
    RECT 498.640 4.600 500.480 1048.040 ;
    RECT 502.320 4.600 504.160 1048.040 ;
    RECT 506.000 4.600 507.840 1048.040 ;
    RECT 509.680 4.600 511.520 1048.040 ;
    RECT 513.360 4.600 515.200 1048.040 ;
    RECT 517.040 4.600 518.880 1048.040 ;
    RECT 520.720 4.600 522.560 1048.040 ;
    RECT 524.400 4.600 526.240 1048.040 ;
    RECT 528.080 4.600 529.920 1048.040 ;
    RECT 531.760 4.600 533.600 1048.040 ;
    RECT 535.440 4.600 537.280 1048.040 ;
    RECT 539.120 4.600 540.960 1048.040 ;
    RECT 542.800 4.600 544.640 1048.040 ;
    RECT 546.480 4.600 548.320 1048.040 ;
    RECT 550.160 4.600 552.000 1048.040 ;
    RECT 553.840 4.600 555.680 1048.040 ;
    RECT 557.520 4.600 559.360 1048.040 ;
    RECT 561.200 4.600 563.040 1048.040 ;
    RECT 564.880 4.600 566.720 1048.040 ;
    RECT 568.560 4.600 570.400 1048.040 ;
    RECT 572.240 4.600 574.080 1048.040 ;
    RECT 575.920 4.600 577.760 1048.040 ;
    RECT 579.600 4.600 581.440 1048.040 ;
    RECT 583.280 4.600 585.120 1048.040 ;
    RECT 586.960 4.600 588.800 1048.040 ;
    RECT 590.640 4.600 592.480 1048.040 ;
    RECT 594.320 4.600 596.160 1048.040 ;
    RECT 598.000 4.600 599.840 1048.040 ;
    RECT 601.680 4.600 603.520 1048.040 ;
    RECT 605.360 4.600 607.200 1048.040 ;
    RECT 609.040 4.600 610.880 1048.040 ;
    RECT 612.720 4.600 614.560 1048.040 ;
    RECT 616.400 4.600 618.240 1048.040 ;
    RECT 620.080 4.600 621.920 1048.040 ;
    RECT 623.760 4.600 625.600 1048.040 ;
    RECT 627.440 4.600 629.280 1048.040 ;
    RECT 631.120 4.600 632.960 1048.040 ;
    RECT 634.800 4.600 636.640 1048.040 ;
    RECT 638.480 4.600 640.320 1048.040 ;
    RECT 642.160 4.600 644.000 1048.040 ;
    RECT 645.840 4.600 647.680 1048.040 ;
    RECT 649.520 4.600 651.360 1048.040 ;
    RECT 653.200 4.600 655.040 1048.040 ;
    RECT 656.880 4.600 658.720 1048.040 ;
    RECT 660.560 4.600 662.400 1048.040 ;
    RECT 664.240 4.600 666.080 1048.040 ;
    RECT 667.920 4.600 669.760 1048.040 ;
    RECT 671.600 4.600 673.440 1048.040 ;
    RECT 675.280 4.600 677.120 1048.040 ;
    RECT 678.960 4.600 680.800 1048.040 ;
    RECT 682.640 4.600 684.480 1048.040 ;
    RECT 686.320 4.600 688.160 1048.040 ;
    RECT 690.000 4.600 691.840 1048.040 ;
    RECT 693.680 4.600 695.520 1048.040 ;
    RECT 697.360 4.600 699.200 1048.040 ;
    RECT 701.040 4.600 702.880 1048.040 ;
    RECT 704.720 4.600 706.560 1048.040 ;
    RECT 708.400 4.600 710.240 1048.040 ;
    RECT 712.080 4.600 713.920 1048.040 ;
    RECT 715.760 4.600 717.600 1048.040 ;
    RECT 719.440 4.600 721.280 1048.040 ;
    RECT 723.120 4.600 724.960 1048.040 ;
    RECT 726.800 4.600 728.640 1048.040 ;
    RECT 730.480 4.600 732.320 1048.040 ;
    RECT 734.160 4.600 736.000 1048.040 ;
    RECT 737.840 4.600 739.680 1048.040 ;
    RECT 741.520 4.600 743.360 1048.040 ;
    RECT 745.200 4.600 747.040 1048.040 ;
    RECT 748.880 4.600 750.720 1048.040 ;
    RECT 752.560 4.600 754.400 1048.040 ;
    RECT 756.240 4.600 758.080 1048.040 ;
    RECT 759.920 4.600 761.760 1048.040 ;
    RECT 763.600 4.600 765.440 1048.040 ;
    RECT 767.280 4.600 769.120 1048.040 ;
    RECT 770.960 4.600 772.800 1048.040 ;
    RECT 774.640 4.600 776.480 1048.040 ;
    RECT 778.320 4.600 780.160 1048.040 ;
    RECT 782.000 4.600 783.840 1048.040 ;
    RECT 785.680 4.600 787.520 1048.040 ;
    RECT 789.360 4.600 791.200 1048.040 ;
    RECT 793.040 4.600 794.880 1048.040 ;
    RECT 796.720 4.600 798.560 1048.040 ;
    RECT 800.400 4.600 802.240 1048.040 ;
    RECT 804.080 4.600 805.920 1048.040 ;
    RECT 807.760 4.600 809.600 1048.040 ;
    RECT 811.440 4.600 813.280 1048.040 ;
    RECT 815.120 4.600 816.960 1048.040 ;
    RECT 818.800 4.600 820.640 1048.040 ;
    RECT 822.480 4.600 824.320 1048.040 ;
    RECT 826.160 4.600 828.000 1048.040 ;
    RECT 829.840 4.600 834.440 1048.040 ;
    LAYER OVERLAP ;
    RECT 0 0 834.440 1052.640 ;
  END
END fakeram130_256x512

END LIBRARY
